//
// Verilog Module mopshub_lib.elink_proc_out_direct
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 18:59:12 09/29/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module elink_proc_out_direct ;


// ### Please start your Verilog code here ### 

endmodule
