//
// Verilog Module mopshub_lib.tb_EPROC_OUT
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 17:17:22 03/16/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
//the test bench should send 8 bits of data with the clock bitCLKx4 
//the data is assigned with a code of 2 bits [00"data, 01"eop, 10"sop, 11"comma]
// dataINrdy is enabled each time the data is available

module tb_EPROC_OUT ;
   // Port Declarations
   wire [1:0] EDATA_OUT;
   wire getDataTrig;
   
    reg [9:0] edataIN; // 10 bits input code+data
    reg dataINrdy;
   
    reg   rst; 
    reg   clk40;     //bitCLK to send the 2bits EdataOUT [clk_40 MB/s]
    reg   clk160;  //bitCLKx4 for 8b/10b encoding [clk_160 MB/s]
    
    reg   swap_output; //No swap equal to 0
    reg   reverse_tx; //normally it is equal to 0 (//LSB send first ) 
    
    wire [1:0] edata_out_s;

// Instances 
assign edata_out_s = U_0.edata_out_s;  
//assign byte= U_0.byte;

EPROC_OUT U_0( 
               .DATA_IN       (edataIN), 
               .DATA_RDY    (dataINrdy),
               .getDataTrig   (getDataTrig), 
               .EDATA_OUT      (EDATA_OUT), 
               .rst           (rst), 
               .bitCLK        (clk40),
               .bitCLKx4      (clk160),
               .swap_outbits  (swap_output),
               .fhCR_REVERSE_10B(reverse_tx)
                ); 
                
  initial begin 
    clk40=0; 
    forever #20 clk40=~clk40; 
  end
  
  initial begin 
    clk160=0; 
    forever #10 clk160=~clk160; 
  end 
  
  
  initial 
  begin
  clk40=1'b1;
  rst = 1'b1;
  #1 rst=!rst;
  
  reverse_tx = 0;
  swap_output  = 0;
  
  edataIN=8'b00010101; 
  dataINrdy=1'b0; 
end
always @(posedge clk40) 
  begin
   $monitor("Time %g   edataIN %b EDATA_OUT %b ",$time, edataIN, EDATA_OUT);
      #2;
      dataINrdy<=1'b1;
      edataIN<=edataIN+1;
      
   end
endmodule
