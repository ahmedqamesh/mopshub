//
// Verilog Module mopshub_lib.Elink_to_FIFO
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 18:57:46 04/02/21
//
// using Mentor Graphics HDL Designer(TM) 2018.1 (Build 12)
//

`resetall
`timescale 1ns/10ps
module Elink_to_FIFO ;


// ### Please start your Verilog code here ### 

endmodule
