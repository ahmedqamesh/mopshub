//
// Verilog Module mopshub_lib.tb_EPROC_OUT_ENC8b10b
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 16:34:52 03/18/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module tb_EPROC_OUT_ENC8b10b ;
  // Port Declarations
  reg   rst; 
  reg   wr_clk;     //bitCLK to send the 2bits EdataOUT [clk_40 MB/s]
  reg   DATA_RDY;
  //EPROC OUT ENC8b10b Signals
  wire [1:0] ENC_EDATA_OUT_2bit;
  wire getDataTrig;
  reg [9:0] GEN_EDATA_10bit; // 10 bits input code+data
  
  //GBTX Emulator
  wire [7:0]  DEC_EDATA_OUT_8bit;
  wire [9:0]  ENC_EDATA_OUT_10bit;
  wire        ko;
  wire        code_err;
  wire        disp_err;
  
  //Data generator Signals
  reg         gen_clk;
  wire        done; 
  wire        wen;
  wire [17:0] GEN_EDATA_18bit;
  

  
  
  data_generator DataGEN(
  .clk_usr  (gen_clk),
  .enable   (~rst),
  .loop_en  (~rst),
  .done     (done),
  .tx_fifo_pfull(1'b0),
  .dout     (GEN_EDATA_18bit),
  .wen      (wen)
  );
  
  
  EPROC_OUT_ENC8b10b U_0( 
  .edataIN       (GEN_EDATA_10bit), 
  .DATA_RDY      (DATA_RDY), //one? CLKx4 after inp_request_trig_out
  .getDataTrig   (getDataTrig), 
  .EDATA_OUT     (ENC_EDATA_OUT_2bit), 
  .rst           (rst), 
  .bitCLK        (wr_clk),  // runs the counters as a normal FIFO clk
  .swap_outbits  (1'b0), //No swap equal to 0
  .fhCR_REVERSE_10B(1'b0)//normally it is equal to 0 (//LSB send first ) enc10bit_r = enc10bit
  ); 
  
  
  GBTX_Emulator U_1( 
  .ko               (ko), 
  .code_err         (code_err), 
  .disp_err         (disp_err), 
  .dataout          (DEC_EDATA_OUT_8bit), 
  .rst              (rst), 
  .datain_valid     (~rst),
  .bitCLK           (wr_clk),
  .enc10bit_out_sig (ENC_EDATA_OUT_10bit),
  .EDATA_2bit       (ENC_EDATA_OUT_2bit),
  .data_10b_in      (10'b0), 
  .data_10b_en      (1'b0)
  );
  
  // clocks           
  initial begin 
    wr_clk=0; 
    forever #1 wr_clk=~wr_clk;
  end
  
  //Generator clk
  initial begin 
    gen_clk=0; 
    forever #4 gen_clk=~gen_clk; 
  end
  
  //Initialization
  initial 
  begin
    DATA_RDY = 1'b0;
    rst = 1'b1;
    #10 rst=!rst;
  end
  
  //initial 
  always@(GEN_EDATA_18bit)
  begin

    #5;
    DATA_RDY = 1'b1;
    GEN_EDATA_10bit = {GEN_EDATA_18bit[17:16],GEN_EDATA_18bit[15:8]};
    #4;//wait 4 wr_clks
    DATA_RDY = 1'b0;
    
    #5;
    GEN_EDATA_10bit = {GEN_EDATA_18bit[17:16],GEN_EDATA_18bit[7:0]};
    DATA_RDY = 1'b1;
    #4;//wait 4 wr_clks
    DATA_RDY = 1'b0;
  end  
endmodule
