`resetall
`timescale 1ns/10ps
module node_readdata_select(
   input   wire    [31:0]  can_rec, 
   input   wire    [31:0] readdata_counter,
   input   wire    [15:0]  readdata0, 
   input   wire    [15:0]  readdata1, 
   input   wire    [15:0]  readdata2, 
   input   wire    [15:0]  readdata3, 
   input   wire    [15:0]  readdata4, 
   input   wire    [15:0]  readdata5, 
   input   wire    [15:0]  readdata6, 
   input   wire    [15:0]  readdata7, 
   input   wire    [15:0]  readdata8, 
   input   wire    [15:0]  readdata9, 
   input   wire    [15:0]  readdata10, 
   input   wire    [15:0]  readdata11, 
   input   wire    [15:0]  readdata12, 
   input   wire    [15:0]  readdata13, 
   input   wire    [15:0]  readdata14, 
   input   wire    [15:0]  readdata15, 
   input   wire    [15:0]  readdata16, 
   input   wire    [15:0]  readdata17, 
   input   wire    [15:0]  readdata18, 
   input   wire    [15:0]  readdata19, 
   input   wire    [15:0]  readdata20, 
   input   wire    [15:0]  readdata21, 
   input   wire    [15:0]  readdata22, 
   input   wire    [15:0]  readdata23, 
   input   wire    [15:0]  readdata24, 
   input   wire    [15:0]  readdata25, 
   input   wire    [15:0]  readdata26, 
   input   wire    [15:0]  readdata27, 
   input   wire    [15:0]  readdata28, 
   input   wire    [15:0]  readdata29, 
   input   wire    [15:0]  readdata30, 
   input   wire    [15:0]  readdata31, 
   
   output   wire   [4:0]  bus_rec_select, 
   output  wire    [15:0]  readdata
);
reg [15:0] readdata_reg ;
reg [15:0] bus_rec_select_reg ;

assign bus_rec_select = bus_rec_select_reg;
assign readdata = readdata_reg;

always @(*)
begin 
 case (readdata_counter)
  31'b01 :
  begin 
    readdata_reg = readdata0;
    bus_rec_select_reg= 5'b00000; 
  end
  31'b010 :
  begin 
    readdata_reg = readdata1;
    bus_rec_select_reg= 5'b00001;
  end
  31'b0100 :
  begin 
    readdata_reg = readdata2;
    bus_rec_select_reg= 5'b00010;
  end
   default : 
   begin 
    readdata_reg = readdata0;
    bus_rec_select_reg= 5'b00000;
  end   
 endcase
end
endmodule
