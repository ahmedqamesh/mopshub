`resetall
`timescale 1ns/10ps
module node_readdata_select( 
   output  wire    [4:0]  can_rec_counter, 
   input   wire    [31:0]  readdata_counter
);

// Internal Declarations
reg [4:0] can_rec_counter_reg ;
assign can_rec_counter = can_rec_counter_reg;

always @(*)
begin 
 case (readdata_counter)
   32'b1: can_rec_counter_reg = 5'h0;
   32'b10: can_rec_counter_reg = 5'h1;
   32'b100: can_rec_counter_reg = 5'h2;
   32'b1000: can_rec_counter_reg = 5'h3;
   32'b10000: can_rec_counter_reg = 5'h4;
   32'b100000: can_rec_counter_reg = 5'h5;
   32'b1000000: can_rec_counter_reg = 5'h6;
   32'b10000000: can_rec_counter_reg = 5'h7;
   32'b100000000: can_rec_counter_reg = 5'h8;
   32'b1000000000: can_rec_counter_reg = 5'h9;
   32'b10000000000: can_rec_counter_reg = 5'hA;
   32'b100000000000: can_rec_counter_reg = 5'hB;
   32'b1000000000000: can_rec_counter_reg = 5'hC;
   32'b10000000000000: can_rec_counter_reg = 5'hD;
   32'b100000000000000: can_rec_counter_reg = 5'hE;
   32'b1000000000000000: can_rec_counter_reg = 5'hF;
   32'b10000000000000000: can_rec_counter_reg = 5'h10;
   32'b100000000000000000: can_rec_counter_reg = 5'h11;
   32'b1000000000000000000: can_rec_counter_reg = 5'h12;
   32'b10000000000000000000: can_rec_counter_reg = 5'h13;
   32'b100000000000000000000: can_rec_counter_reg = 5'h14;
   32'b1000000000000000000000: can_rec_counter_reg = 5'h15;
   32'b10000000000000000000000: can_rec_counter_reg = 5'h16;
   32'b100000000000000000000000: can_rec_counter_reg = 5'h17;
   32'b1000000000000000000000000: can_rec_counter_reg = 5'h18;
   32'b10000000000000000000000000: can_rec_counter_reg = 5'h19;
   32'b100000000000000000000000000: can_rec_counter_reg = 5'h1A;
   32'b1000000000000000000000000000: can_rec_counter_reg = 5'h1B;
   32'b10000000000000000000000000000: can_rec_counter_reg = 5'h1C;
   32'b100000000000000000000000000000: can_rec_counter_reg = 5'h1D;
   32'b1000000000000000000000000000000: can_rec_counter_reg = 5'h1E;
   32'b10000000000000000000000000000000: can_rec_counter_reg = 5'h1F;
   endcase   
end
endmodule
