//
// Verilog Module mopshub_lib.demux_1_8_8bit
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 13:38:43 06/14/23
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module demux_1_8_8bit ;


// ### Please start your Verilog code here ### 

endmodule
