//
// Verilog Module mopshub_lib.tb_ring_counter
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 13:08:45 01/13/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module tb_readdata_counter;
	// Inputs
	reg clock;
	reg reset;
	// Outputs
  wire[31:0] readdata_counter;
	// Instantiate the Unit Under Test (UUT)
	node_readdata_counter uut (
      .clock(clock), 
      .reset(reset), 
      .readdata_counter(readdata_counter)
	);
 always #1 clock = ~clock;
	initial begin
	  $monitor($time, " clock=%1b,reset=%1b,readdata_counter=%b",clock,reset,readdata_counter);
		// Initialize Inputs
    clock = 0;  
	  reset = 0;
 
	#1 reset = 1;
	#1 reset = 0; 
	
    end  
    
endmodule
