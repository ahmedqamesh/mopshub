//
// Verilog Module mopshub_lib.tb_fifo_to_2K_18bit_wide
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 13:52:37 03/01/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module tb_fifo_to_2K_18bit_wide ;
  
  parameter DATA_WIDTH=18;
  parameter ADDRESS_WIDTH = 11;
  parameter FIFO_DEPTH = 16 ;//(1 << ADDRESS_WIDTH);// the FIFO depth is  2K (2^11)

  wire [DATA_WIDTH-1:0] dout;
  wire almost_full,full,empty;
  
  
  reg [DATA_WIDTH-1:0] din;
  reg rd_en,wr_en,rd_clk,wr_clk;
  reg rst;
  
  wire [3:0] r_ptr,w_ptr,ptr_diff;
  
  assign r_ptr=fifo2K_18bit_wide.r_ptr;
  assign w_ptr=fifo2K_18bit_wide.w_ptr;
  assign ptr_diff=fifo2K_18bit_wide.ptr_diff;
  assign r_next_en=fifo2K_18bit_wide.r_next_en;
  assign w_next_en=fifo2K_18bit_wide.w_next_en;

  
  fh_epath_fifo2K_18bit_wide fifo2K_18bit_wide(dout,full,empty,
  
  almost_full,din,rd_en,wr_en,rd_clk,wr_clk,rst);
  
  
  
  
  //initial #5000 $stop;
  initial begin 
    #10 rd_clk=0; 
    forever #10 rd_clk=~rd_clk; 
  end
  
  initial begin 
    #5 wr_clk=0; 
    forever #50 wr_clk=~wr_clk; 
  end  
  
  initial begin din=1;
  @(posedge wr_en);
    repeat(20) @(posedge wr_clk) din=din+2;
    repeat(20) @(posedge wr_clk) din=din-1;
    end
  
  initial begin rst=1;#30 rst=0;end 
  initial begin fork #50 wr_en=1; #1800 wr_en=0; #2500 wr_en=1 ; join end            
  initial begin
    $monitor("din %d dout %d",din,dout);
    fork #50 rd_en=0; 
    #1850 rd_en=1; 
    #2400 rd_en=0; 
    #2500 rd_en=1; 
  join end
                
endmodule