`resetall
`timescale 1ns/10ps
module tb_readdata_select;
	// Inputs
	 reg clock;
	 reg reset;
	
	// Outputs
   wire   [4:0]  can_rec_counter;
	// Instantiate the Unit Under Test (UUT)
	test_block uut (
      .can_rec_counter(can_rec_counter),                                     
      .clock(clock), 
      .reset(reset) 
	);
	always #1 clock = ~clock;
  initial begin
    $monitor($time,  " : clock= %g reset = %b can_rec_counter = %d",
              clock,reset, can_rec_counter);
		// Initialize Inputs
    clock = 0;  
	#1 reset = 1;
	#1 reset = 0; 
  end 
endmodule
