//
// Verilog Module mopshub_lib.data_gen_elink_SM
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 18:41:35 06/21/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module data_gen_elink_SM ;


// ### Please start your Verilog code here ### 

endmodule
