//
// Verilog Module mopshub_lib.data_gen_elink
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 19:02:34 06/21/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module data_gen_elink ;


// ### Please start your Verilog code here ### 

endmodule
