--! This file is part of the FELIX firmware distribution (https://gitlab.cern.ch/atlas-tdaq-felix/firmware/).
--! Copyright (C) 2001-2021 CERN for the benefit of the ATLAS collaboration.
--! Authors:
--!               Mark Donszelmann
--!               Andrea Borga
--!               Soo Ryu
--!               Kai Chen
--!               Israel Grayzman
--!               Rene Habraken
--!               Alexander Paramonov
--!               RHabraken
--!               Nayib Boukadida
--!               Alessandra Camplani
--!               Elena Zhivun
--!               Mesfin Gebyehu
--!               Rene
--!               Thei Wijnen
--!               Ohad Shaked
--!               Alessandro Thea
--!               mtrovato
--!               Frans Schreuder
--! 
--!   Licensed under the Apache License, Version 2.0 (the "License");
--!   you may not use this file except in compliance with the License.
--!   You may obtain a copy of the License at
--!
--!       http://www.apache.org/licenses/LICENSE-2.0
--!
--!   Unless required by applicable law or agreed to in writing, software
--!   distributed under the License is distributed on an "AS IS" BASIS,
--!   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--!   See the License for the specific language governing permissions and
--!   limitations under the License.
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- DO NOT EDIT THIS FILE
-- 
-- This file was generated from template '../../../sources/templates/jinja/pcie_package.vhd.template'
-- and register map ../../../sources/templates/yaml/registers-5.0.yaml, version 5.0
-- by the script 'wuppercodegen', version: 0.8.6,
-- using the following commandline:
-- 
-- ../../../WupperCodeGen/wuppercodegen/cli.py ../../../sources/templates/yaml/registers-5.0.yaml ../../../sources/templates/jinja/pcie_package.vhd.template ../../../sources/templates/generated/pcie_package.vhd
-- 
-- Please do NOT edit this file, but edit the source file at '../../../sources/templates/jinja/pcie_package.vhd.template'
-- 
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************


--!------------------------------------------------------------------------------
--!
--!           NIKHEF - National Institute for Subatomic Physics
--!
--!                       Electronics Department
--!
--!-----------------------------------------------------------------------------
--! @class pcie_package
--!
--!
--! @author      Andrea Borga    (andrea.borga@nikhef.nl)<br>
--!              Frans Schreuder (frans.schreuder@nikhef.nl)
--!
--!
--! @date        07/01/2015    created
--!
--! @version     1.0
--!
--! @brief
--! This package contains the data types for the PCIe DMA core, as well as some
--! constants, addresses and register types for the application.
--!
--!
--! @detail
--!
--!-----------------------------------------------------------------------------
--! @TODO
--!
--!
--! ------------------------------------------------------------------------------
--!

--! @brief ieee



library ieee;
use ieee.numeric_std.all;
--use ieee.std_logic_unsigned.all;
use ieee.std_logic_1164.all;

use work.centralRouter_package.all;
use work.data_width_package.all;

package pcie_package is

  function to_sl( A: std_logic_vector) return std_logic ;
  function or_reduce(slv : in std_logic_vector) return std_logic ;
  --
  -- PCIe DMA core: AXI-4 Stream interface
  type axis_type is record
    tdata   : std_logic_vector(PCIE_DATA_WIDTH-1 downto 0);
    tkeep   : std_logic_vector(15 downto 0);
    tuser   : std_logic_vector(182 downto 0);
    tlast   : std_logic;
    tvalid  : std_logic;
    state   : std_logic_vector(2 downto 0); --debugging purposes, connected to ILA
  end record;

  type axis_r_type is record
    tready: std_logic;
  end record;

  --
  -- PCIe DMA core: descriptors
  type dma_descriptor_type is record
    start_address   : std_logic_vector(63 downto 0);
    end_address     : std_logic_vector(63 downto 0);
    dword_count     : std_logic_vector(10 downto 0);
    read_not_write  : std_logic;     --1 means this is a read descriptor, 0: write descriptor
    enable          : std_logic;     --descriptor is valid
    wrap_around     : std_logic;     --1 means when end is reached, keep enabled and start over
    evencycle_pc    : std_logic;     --For every time the pc pointer overflows, this bit toggles.
    pc_pointer      : std_logic_vector(63 downto 0); --Last address that the PC has read / written. For write: overflow and read until this cycle.
    pc_pointer_updated : std_logic;  --Pulse when the pc_pointer is written
  end record;

  type dma_descriptors_type is array (natural range <>) of dma_descriptor_type;

  type dma_status_type is record
    current_address : std_logic_vector(63 downto 0);
    evencycle_dma   : std_logic;     --For every time the current_address overflows, this bit toggles
    address_wrapped : std_logic;
  end record;

  type dma_statuses_type is array(natural range <>) of dma_status_type;

  --
  -- PCIe DMA core: Interrupt Vectors
  type interrupt_vector_type is record
    int_vec_add  : std_logic_vector(63 downto 0);
    int_vec_data : std_logic_vector(31 downto 0);
    int_vec_ctrl : std_logic_vector(31 downto 0);
  end record;

  type interrupt_vectors_type is array (natural range <>) of interrupt_vector_type;
  
  type slv_array is array (natural range <>) of std_logic_vector(PCIE_DATA_WIDTH-1 downto 0);
  type slv12_array is array (natural range <>) of std_logic_vector(11 downto 0);

  --! Address Offset assignment
  --! --> BAR0 User Application Registers Addresses
  -- ### BAR0 registers: start
  constant REG_DESCRIPTOR_0        : std_logic_vector(19 downto 0) := x"00000";
  constant REG_DESCRIPTOR_0a       : std_logic_vector(19 downto 0) := x"00010";
  constant REG_DESCRIPTOR_1        : std_logic_vector(19 downto 0) := x"00020";
  constant REG_DESCRIPTOR_1a       : std_logic_vector(19 downto 0) := x"00030";
  constant REG_DESCRIPTOR_2        : std_logic_vector(19 downto 0) := x"00040";
  constant REG_DESCRIPTOR_2a       : std_logic_vector(19 downto 0) := x"00050";
  constant REG_DESCRIPTOR_3        : std_logic_vector(19 downto 0) := x"00060";
  constant REG_DESCRIPTOR_3a       : std_logic_vector(19 downto 0) := x"00070";
  constant REG_DESCRIPTOR_4        : std_logic_vector(19 downto 0) := x"00080";
  constant REG_DESCRIPTOR_4a       : std_logic_vector(19 downto 0) := x"00090";
  constant REG_DESCRIPTOR_5        : std_logic_vector(19 downto 0) := x"000A0";
  constant REG_DESCRIPTOR_5a       : std_logic_vector(19 downto 0) := x"000B0";
  constant REG_DESCRIPTOR_6        : std_logic_vector(19 downto 0) := x"000C0";
  constant REG_DESCRIPTOR_6a       : std_logic_vector(19 downto 0) := x"000D0";
  constant REG_DESCRIPTOR_7        : std_logic_vector(19 downto 0) := x"000E0";
  constant REG_DESCRIPTOR_7a       : std_logic_vector(19 downto 0) := x"000F0";
  constant REG_DESCRIPTOR_8        : std_logic_vector(19 downto 0) := x"00100";
  constant REG_DESCRIPTOR_8a       : std_logic_vector(19 downto 0) := x"00110";
  constant REG_DESCRIPTOR_9        : std_logic_vector(19 downto 0) := x"00120";
  constant REG_DESCRIPTOR_9a       : std_logic_vector(19 downto 0) := x"00130";
  constant REG_DESCRIPTOR_10       : std_logic_vector(19 downto 0) := x"00140";
  constant REG_DESCRIPTOR_10a      : std_logic_vector(19 downto 0) := x"00150";
  constant REG_DESCRIPTOR_11       : std_logic_vector(19 downto 0) := x"00160";
  constant REG_DESCRIPTOR_11a      : std_logic_vector(19 downto 0) := x"00170";
  constant REG_DESCRIPTOR_12       : std_logic_vector(19 downto 0) := x"00180";
  constant REG_DESCRIPTOR_12a      : std_logic_vector(19 downto 0) := x"00190";
  constant REG_DESCRIPTOR_13       : std_logic_vector(19 downto 0) := x"001A0";
  constant REG_DESCRIPTOR_13a      : std_logic_vector(19 downto 0) := x"001B0";
  constant REG_DESCRIPTOR_14       : std_logic_vector(19 downto 0) := x"001C0";
  constant REG_DESCRIPTOR_14a      : std_logic_vector(19 downto 0) := x"001D0";
  constant REG_DESCRIPTOR_15       : std_logic_vector(19 downto 0) := x"001E0";
  constant REG_DESCRIPTOR_15a      : std_logic_vector(19 downto 0) := x"001F0";
  constant REG_STATUS_0            : std_logic_vector(19 downto 0) := x"00200";
  constant REG_STATUS_1            : std_logic_vector(19 downto 0) := x"00210";
  constant REG_STATUS_2            : std_logic_vector(19 downto 0) := x"00220";
  constant REG_STATUS_3            : std_logic_vector(19 downto 0) := x"00230";
  constant REG_STATUS_4            : std_logic_vector(19 downto 0) := x"00240";
  constant REG_STATUS_5            : std_logic_vector(19 downto 0) := x"00250";
  constant REG_STATUS_6            : std_logic_vector(19 downto 0) := x"00260";
  constant REG_STATUS_7            : std_logic_vector(19 downto 0) := x"00270";
  constant REG_STATUS_8            : std_logic_vector(19 downto 0) := x"00280";
  constant REG_STATUS_9            : std_logic_vector(19 downto 0) := x"00290";
  constant REG_STATUS_10           : std_logic_vector(19 downto 0) := x"002A0";
  constant REG_STATUS_11           : std_logic_vector(19 downto 0) := x"002B0";
  constant REG_STATUS_12           : std_logic_vector(19 downto 0) := x"002C0";
  constant REG_STATUS_13           : std_logic_vector(19 downto 0) := x"002D0";
  constant REG_STATUS_14           : std_logic_vector(19 downto 0) := x"002E0";
  constant REG_STATUS_15           : std_logic_vector(19 downto 0) := x"002F0";
  constant REG_BAR0                : std_logic_vector(19 downto 0) := x"00300";
  constant REG_BAR1                : std_logic_vector(19 downto 0) := x"00310";
  constant REG_BAR2                : std_logic_vector(19 downto 0) := x"00320";
  constant REG_DESCRIPTOR_ENABLE   : std_logic_vector(19 downto 0) := x"00400";
  constant REG_FIFO_FLUSH          : std_logic_vector(19 downto 0) := x"00410";
  constant REG_DMA_RESET           : std_logic_vector(19 downto 0) := x"00420";
  constant REG_SOFT_RESET          : std_logic_vector(19 downto 0) := x"00430";
  constant REG_REGISTER_RESET      : std_logic_vector(19 downto 0) := x"00440";
  constant REG_FROMHOST_FULL_THRESH: std_logic_vector(19 downto 0) := x"00450";
  constant REG_TOHOST_FULL_THRESH  : std_logic_vector(19 downto 0) := x"00460";
  constant REG_BUSY_THRESH_ASSERT  : std_logic_vector(19 downto 0) := x"00470";
  constant REG_BUSY_THRESH_NEGATE  : std_logic_vector(19 downto 0) := x"00480";
  constant REG_BUSY_STATUS         : std_logic_vector(19 downto 0) := x"00490";
  constant REG_PC_PTR_GAP          : std_logic_vector(19 downto 0) := x"004A0";
  
  -- BAR0 registers: end

  --! Address Offset assignment
  --! --> BAR1 User Application Registers Addresses
  -- ### BAR1 registers: start
     -- interrupt vectors
  constant REG_INT_VEC_00          : std_logic_vector(19 downto 0) := x"00000";
  constant REG_INT_VEC_01          : std_logic_vector(19 downto 0) := x"00010";
  constant REG_INT_VEC_02          : std_logic_vector(19 downto 0) := x"00020";
  constant REG_INT_VEC_03          : std_logic_vector(19 downto 0) := x"00030";
  constant REG_INT_VEC_04          : std_logic_vector(19 downto 0) := x"00040";
  constant REG_INT_VEC_05          : std_logic_vector(19 downto 0) := x"00050";
  constant REG_INT_VEC_06          : std_logic_vector(19 downto 0) := x"00060";
  constant REG_INT_VEC_07          : std_logic_vector(19 downto 0) := x"00070";
  constant REG_INT_VEC_08          : std_logic_vector(19 downto 0) := x"00080";
  constant REG_INT_VEC_09          : std_logic_vector(19 downto 0) := x"00090";
  constant REG_INT_VEC_10          : std_logic_vector(19 downto 0) := x"000A0";
  constant REG_INT_VEC_11          : std_logic_vector(19 downto 0) := x"000B0";
  constant REG_INT_VEC_12          : std_logic_vector(19 downto 0) := x"000C0";
  constant REG_INT_VEC_13          : std_logic_vector(19 downto 0) := x"000D0";
  constant REG_INT_VEC_14          : std_logic_vector(19 downto 0) := x"000E0";
  constant REG_INT_VEC_15          : std_logic_vector(19 downto 0) := x"000F0";
  constant REG_INT_TAB_EN          : std_logic_vector(19 downto 0) := x"00100";
  -- BAR1 registers: end


  --! Address Offset assignment
  --! --> BAR2 User Application Registers Addresses
  --! -- leave 16x8 = 128 bits space per register
  ------------------------------------
  ---- ## GENERATED code BEGIN #1 ----
  ------------------------------------

  --** Bar2

  --** GenericBoardInformation
  constant REG_REG_MAP_VERSION                : std_logic_vector(19 downto 0) := x"00000";
  constant REG_BOARD_ID_TIMESTAMP             : std_logic_vector(19 downto 0) := x"00010";
  constant REG_GIT_COMMIT_TIME                : std_logic_vector(19 downto 0) := x"00030";
  constant REG_GIT_TAG                        : std_logic_vector(19 downto 0) := x"00040";
  constant REG_GIT_COMMIT_NUMBER              : std_logic_vector(19 downto 0) := x"00050";
  constant REG_GIT_HASH                       : std_logic_vector(19 downto 0) := x"00060";
  constant REG_STATUS_LEDS                    : std_logic_vector(19 downto 0) := x"00070";
  constant REG_GENERIC_CONSTANTS              : std_logic_vector(19 downto 0) := x"00080";
  constant REG_NUM_OF_CHANNELS                : std_logic_vector(19 downto 0) := x"00090";
  constant REG_CARD_TYPE                      : std_logic_vector(19 downto 0) := x"000a0";
  constant REG_GENERATE_GBT                   : std_logic_vector(19 downto 0) := x"000c0";
  constant REG_OPTO_TRX_NUM                   : std_logic_vector(19 downto 0) := x"000d0";
  constant REG_GENERATE_TTC_EMU               : std_logic_vector(19 downto 0) := x"000e0";

  --** INCLUDE_EGROUPS
  constant REG_INCLUDE_EGROUP_0               : std_logic_vector(19 downto 0) := x"00100";
  constant REG_INCLUDE_EGROUP_1               : std_logic_vector(19 downto 0) := x"00110";
  constant REG_INCLUDE_EGROUP_2               : std_logic_vector(19 downto 0) := x"00120";
  constant REG_INCLUDE_EGROUP_3               : std_logic_vector(19 downto 0) := x"00130";
  constant REG_INCLUDE_EGROUP_4               : std_logic_vector(19 downto 0) := x"00140";
  constant REG_INCLUDE_EGROUP_5               : std_logic_vector(19 downto 0) := x"00150";
  constant REG_INCLUDE_EGROUP_6               : std_logic_vector(19 downto 0) := x"00160";
  constant REG_WIDE_MODE                      : std_logic_vector(19 downto 0) := x"00170";
  constant REG_FIRMWARE_MODE                  : std_logic_vector(19 downto 0) := x"00190";
  constant REG_GTREFCLK_SOURCE                : std_logic_vector(19 downto 0) := x"001a0";
  constant REG_CR_GENERICS                    : std_logic_vector(19 downto 0) := x"001b0";
  constant REG_BLOCKSIZE                      : std_logic_vector(19 downto 0) := x"001c0";
  constant REG_PCIE_ENDPOINT                  : std_logic_vector(19 downto 0) := x"001d0";
  constant REG_CHUNK_TRAILER_32B              : std_logic_vector(19 downto 0) := x"001e0";
  constant REG_NUMBER_OF_PCIE_ENDPOINTS       : std_logic_vector(19 downto 0) := x"001f0";
  constant REG_AXI_STREAMS_TOHOST             : std_logic_vector(19 downto 0) := x"00200";
  constant REG_AXI_STREAMS_FROMHOST           : std_logic_vector(19 downto 0) := x"00210";
  constant REG_FROMHOST_LENGTH_IS_5BIT        : std_logic_vector(19 downto 0) := x"00220";
  constant REG_FULLMODE_HALFRATE              : std_logic_vector(19 downto 0) := x"00230";
  constant REG_SUPPORT_HDLC_DELAY             : std_logic_vector(19 downto 0) := x"00240";

  --** CRToHostControlsAndMonitors
  constant REG_TIMEOUT_CTRL                   : std_logic_vector(19 downto 0) := x"00800";
  constant REG_MAX_TIMEOUT                    : std_logic_vector(19 downto 0) := x"00810";
  constant REG_CRTOHOST_FIFO_STATUS           : std_logic_vector(19 downto 0) := x"00820";
  constant REG_CRTOHOST_DMA_DESCRIPTOR_1      : std_logic_vector(19 downto 0) := x"00830";
  constant REG_CRTOHOST_DMA_DESCRIPTOR_2      : std_logic_vector(19 downto 0) := x"00840";

  --** CRFromHostControlsAndMonitors
  constant REG_CRFROMHOST_FIFO_STATUS         : std_logic_vector(19 downto 0) := x"01000";

  --** BROADCAST_ENABLE_GEN
  constant REG_BROADCAST_ENABLE_00            : std_logic_vector(19 downto 0) := x"01010";
  constant REG_BROADCAST_ENABLE_01            : std_logic_vector(19 downto 0) := x"01020";
  constant REG_BROADCAST_ENABLE_02            : std_logic_vector(19 downto 0) := x"01030";
  constant REG_BROADCAST_ENABLE_03            : std_logic_vector(19 downto 0) := x"01040";
  constant REG_BROADCAST_ENABLE_04            : std_logic_vector(19 downto 0) := x"01050";
  constant REG_BROADCAST_ENABLE_05            : std_logic_vector(19 downto 0) := x"01060";
  constant REG_BROADCAST_ENABLE_06            : std_logic_vector(19 downto 0) := x"01070";
  constant REG_BROADCAST_ENABLE_07            : std_logic_vector(19 downto 0) := x"01080";
  constant REG_BROADCAST_ENABLE_08            : std_logic_vector(19 downto 0) := x"01090";
  constant REG_BROADCAST_ENABLE_09            : std_logic_vector(19 downto 0) := x"010a0";
  constant REG_BROADCAST_ENABLE_10            : std_logic_vector(19 downto 0) := x"010b0";
  constant REG_BROADCAST_ENABLE_11            : std_logic_vector(19 downto 0) := x"010c0";
  constant REG_BROADCAST_ENABLE_12            : std_logic_vector(19 downto 0) := x"010d0";
  constant REG_BROADCAST_ENABLE_13            : std_logic_vector(19 downto 0) := x"010e0";
  constant REG_BROADCAST_ENABLE_14            : std_logic_vector(19 downto 0) := x"010f0";
  constant REG_BROADCAST_ENABLE_15            : std_logic_vector(19 downto 0) := x"01100";
  constant REG_BROADCAST_ENABLE_16            : std_logic_vector(19 downto 0) := x"01110";
  constant REG_BROADCAST_ENABLE_17            : std_logic_vector(19 downto 0) := x"01120";
  constant REG_BROADCAST_ENABLE_18            : std_logic_vector(19 downto 0) := x"01130";
  constant REG_BROADCAST_ENABLE_19            : std_logic_vector(19 downto 0) := x"01140";
  constant REG_BROADCAST_ENABLE_20            : std_logic_vector(19 downto 0) := x"01150";
  constant REG_BROADCAST_ENABLE_21            : std_logic_vector(19 downto 0) := x"01160";
  constant REG_BROADCAST_ENABLE_22            : std_logic_vector(19 downto 0) := x"01170";
  constant REG_BROADCAST_ENABLE_23            : std_logic_vector(19 downto 0) := x"01180";
  constant REG_CRFROMHOST_RESET               : std_logic_vector(19 downto 0) := x"01190";

  --** DecodingControlsAndMonitors

  --** PATH_HAS_STREAM_ID
  constant REG_LINK_00_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02000";
  constant REG_LINK_01_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02010";
  constant REG_LINK_02_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02020";
  constant REG_LINK_03_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02030";
  constant REG_LINK_04_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02040";
  constant REG_LINK_05_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02050";
  constant REG_LINK_06_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02060";
  constant REG_LINK_07_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02070";
  constant REG_LINK_08_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02080";
  constant REG_LINK_09_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02090";
  constant REG_LINK_10_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"020a0";
  constant REG_LINK_11_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"020b0";
  constant REG_LINK_12_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"020c0";
  constant REG_LINK_13_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"020d0";
  constant REG_LINK_14_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"020e0";
  constant REG_LINK_15_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"020f0";
  constant REG_LINK_16_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02100";
  constant REG_LINK_17_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02110";
  constant REG_LINK_18_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02120";
  constant REG_LINK_19_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02130";
  constant REG_LINK_20_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02140";
  constant REG_LINK_21_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02150";
  constant REG_LINK_22_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02160";
  constant REG_LINK_23_HAS_STREAM_ID          : std_logic_vector(19 downto 0) := x"02170";

  --** DECODING_LINK_STATUS_ARR
  constant REG_DECODING_LINK_ALIGNED_00       : std_logic_vector(19 downto 0) := x"02180";
  constant REG_DECODING_LINK_ALIGNED_01       : std_logic_vector(19 downto 0) := x"02190";
  constant REG_DECODING_LINK_ALIGNED_02       : std_logic_vector(19 downto 0) := x"021a0";
  constant REG_DECODING_LINK_ALIGNED_03       : std_logic_vector(19 downto 0) := x"021b0";
  constant REG_DECODING_LINK_ALIGNED_04       : std_logic_vector(19 downto 0) := x"021c0";
  constant REG_DECODING_LINK_ALIGNED_05       : std_logic_vector(19 downto 0) := x"021d0";
  constant REG_DECODING_LINK_ALIGNED_06       : std_logic_vector(19 downto 0) := x"021e0";
  constant REG_DECODING_LINK_ALIGNED_07       : std_logic_vector(19 downto 0) := x"021f0";
  constant REG_DECODING_LINK_ALIGNED_08       : std_logic_vector(19 downto 0) := x"02200";
  constant REG_DECODING_LINK_ALIGNED_09       : std_logic_vector(19 downto 0) := x"02210";
  constant REG_DECODING_LINK_ALIGNED_10       : std_logic_vector(19 downto 0) := x"02220";
  constant REG_DECODING_LINK_ALIGNED_11       : std_logic_vector(19 downto 0) := x"02230";
  constant REG_DECODING_LINK_ALIGNED_12       : std_logic_vector(19 downto 0) := x"02240";
  constant REG_DECODING_LINK_ALIGNED_13       : std_logic_vector(19 downto 0) := x"02250";
  constant REG_DECODING_LINK_ALIGNED_14       : std_logic_vector(19 downto 0) := x"02260";
  constant REG_DECODING_LINK_ALIGNED_15       : std_logic_vector(19 downto 0) := x"02270";
  constant REG_DECODING_LINK_ALIGNED_16       : std_logic_vector(19 downto 0) := x"02280";
  constant REG_DECODING_LINK_ALIGNED_17       : std_logic_vector(19 downto 0) := x"02290";
  constant REG_DECODING_LINK_ALIGNED_18       : std_logic_vector(19 downto 0) := x"022a0";
  constant REG_DECODING_LINK_ALIGNED_19       : std_logic_vector(19 downto 0) := x"022b0";
  constant REG_DECODING_LINK_ALIGNED_20       : std_logic_vector(19 downto 0) := x"022c0";
  constant REG_DECODING_LINK_ALIGNED_21       : std_logic_vector(19 downto 0) := x"022d0";
  constant REG_DECODING_LINK_ALIGNED_22       : std_logic_vector(19 downto 0) := x"022e0";
  constant REG_DECODING_LINK_ALIGNED_23       : std_logic_vector(19 downto 0) := x"022f0";

  --** DECODING_EGROUP_CTRL_GEN

  --** DECODING_EGROUP
  constant REG_DECODING_LINK00_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"02300";
  constant REG_DECODING_LINK00_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"02310";
  constant REG_DECODING_LINK00_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"02320";
  constant REG_DECODING_LINK00_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"02330";
  constant REG_DECODING_LINK00_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"02340";
  constant REG_DECODING_LINK00_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"02350";
  constant REG_DECODING_LINK00_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"02360";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK01_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"02370";
  constant REG_DECODING_LINK01_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"02380";
  constant REG_DECODING_LINK01_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"02390";
  constant REG_DECODING_LINK01_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"023a0";
  constant REG_DECODING_LINK01_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"023b0";
  constant REG_DECODING_LINK01_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"023c0";
  constant REG_DECODING_LINK01_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"023d0";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK02_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"023e0";
  constant REG_DECODING_LINK02_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"023f0";
  constant REG_DECODING_LINK02_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"02400";
  constant REG_DECODING_LINK02_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"02410";
  constant REG_DECODING_LINK02_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"02420";
  constant REG_DECODING_LINK02_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"02430";
  constant REG_DECODING_LINK02_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"02440";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK03_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"02450";
  constant REG_DECODING_LINK03_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"02460";
  constant REG_DECODING_LINK03_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"02470";
  constant REG_DECODING_LINK03_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"02480";
  constant REG_DECODING_LINK03_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"02490";
  constant REG_DECODING_LINK03_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"024a0";
  constant REG_DECODING_LINK03_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"024b0";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK04_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"024c0";
  constant REG_DECODING_LINK04_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"024d0";
  constant REG_DECODING_LINK04_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"024e0";
  constant REG_DECODING_LINK04_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"024f0";
  constant REG_DECODING_LINK04_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"02500";
  constant REG_DECODING_LINK04_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"02510";
  constant REG_DECODING_LINK04_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"02520";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK05_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"02530";
  constant REG_DECODING_LINK05_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"02540";
  constant REG_DECODING_LINK05_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"02550";
  constant REG_DECODING_LINK05_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"02560";
  constant REG_DECODING_LINK05_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"02570";
  constant REG_DECODING_LINK05_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"02580";
  constant REG_DECODING_LINK05_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"02590";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK06_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"025a0";
  constant REG_DECODING_LINK06_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"025b0";
  constant REG_DECODING_LINK06_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"025c0";
  constant REG_DECODING_LINK06_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"025d0";
  constant REG_DECODING_LINK06_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"025e0";
  constant REG_DECODING_LINK06_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"025f0";
  constant REG_DECODING_LINK06_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"02600";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK07_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"02610";
  constant REG_DECODING_LINK07_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"02620";
  constant REG_DECODING_LINK07_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"02630";
  constant REG_DECODING_LINK07_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"02640";
  constant REG_DECODING_LINK07_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"02650";
  constant REG_DECODING_LINK07_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"02660";
  constant REG_DECODING_LINK07_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"02670";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK08_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"02680";
  constant REG_DECODING_LINK08_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"02690";
  constant REG_DECODING_LINK08_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"026a0";
  constant REG_DECODING_LINK08_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"026b0";
  constant REG_DECODING_LINK08_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"026c0";
  constant REG_DECODING_LINK08_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"026d0";
  constant REG_DECODING_LINK08_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"026e0";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK09_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"026f0";
  constant REG_DECODING_LINK09_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"02700";
  constant REG_DECODING_LINK09_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"02710";
  constant REG_DECODING_LINK09_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"02720";
  constant REG_DECODING_LINK09_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"02730";
  constant REG_DECODING_LINK09_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"02740";
  constant REG_DECODING_LINK09_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"02750";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK10_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"02760";
  constant REG_DECODING_LINK10_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"02770";
  constant REG_DECODING_LINK10_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"02780";
  constant REG_DECODING_LINK10_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"02790";
  constant REG_DECODING_LINK10_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"027a0";
  constant REG_DECODING_LINK10_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"027b0";
  constant REG_DECODING_LINK10_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"027c0";

  --** DECODING_EGROUP
  constant REG_DECODING_LINK11_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"027d0";
  constant REG_DECODING_LINK11_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"027e0";
  constant REG_DECODING_LINK11_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"027f0";
  constant REG_DECODING_LINK11_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"02800";
  constant REG_DECODING_LINK11_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"02810";
  constant REG_DECODING_LINK11_EGROUP5_CTRL   : std_logic_vector(19 downto 0) := x"02820";
  constant REG_DECODING_LINK11_EGROUP6_CTRL   : std_logic_vector(19 downto 0) := x"02830";

  --** MINI_EGROUP_TOHOST_GEN
  constant REG_MINI_EGROUP_TOHOST_00          : std_logic_vector(19 downto 0) := x"02840";
  constant REG_MINI_EGROUP_TOHOST_01          : std_logic_vector(19 downto 0) := x"02850";
  constant REG_MINI_EGROUP_TOHOST_02          : std_logic_vector(19 downto 0) := x"02860";
  constant REG_MINI_EGROUP_TOHOST_03          : std_logic_vector(19 downto 0) := x"02870";
  constant REG_MINI_EGROUP_TOHOST_04          : std_logic_vector(19 downto 0) := x"02880";
  constant REG_MINI_EGROUP_TOHOST_05          : std_logic_vector(19 downto 0) := x"02890";
  constant REG_MINI_EGROUP_TOHOST_06          : std_logic_vector(19 downto 0) := x"028a0";
  constant REG_MINI_EGROUP_TOHOST_07          : std_logic_vector(19 downto 0) := x"028b0";
  constant REG_MINI_EGROUP_TOHOST_08          : std_logic_vector(19 downto 0) := x"028c0";
  constant REG_MINI_EGROUP_TOHOST_09          : std_logic_vector(19 downto 0) := x"028d0";
  constant REG_MINI_EGROUP_TOHOST_10          : std_logic_vector(19 downto 0) := x"028e0";
  constant REG_MINI_EGROUP_TOHOST_11          : std_logic_vector(19 downto 0) := x"028f0";
  constant REG_MINI_EGROUP_TOHOST_12          : std_logic_vector(19 downto 0) := x"02900";
  constant REG_MINI_EGROUP_TOHOST_13          : std_logic_vector(19 downto 0) := x"02910";
  constant REG_MINI_EGROUP_TOHOST_14          : std_logic_vector(19 downto 0) := x"02920";
  constant REG_MINI_EGROUP_TOHOST_15          : std_logic_vector(19 downto 0) := x"02930";
  constant REG_MINI_EGROUP_TOHOST_16          : std_logic_vector(19 downto 0) := x"02940";
  constant REG_MINI_EGROUP_TOHOST_17          : std_logic_vector(19 downto 0) := x"02950";
  constant REG_MINI_EGROUP_TOHOST_18          : std_logic_vector(19 downto 0) := x"02960";
  constant REG_MINI_EGROUP_TOHOST_19          : std_logic_vector(19 downto 0) := x"02970";
  constant REG_MINI_EGROUP_TOHOST_20          : std_logic_vector(19 downto 0) := x"02980";
  constant REG_MINI_EGROUP_TOHOST_21          : std_logic_vector(19 downto 0) := x"02990";
  constant REG_MINI_EGROUP_TOHOST_22          : std_logic_vector(19 downto 0) := x"029a0";
  constant REG_MINI_EGROUP_TOHOST_23          : std_logic_vector(19 downto 0) := x"029b0";
  constant REG_TTC_TOHOST_ENABLE              : std_logic_vector(19 downto 0) := x"029c0";
  constant REG_DECODING_REVERSE_10B           : std_logic_vector(19 downto 0) := x"029d0";

  --** YARR_DEBUG_ALLEGROUP_TOHOST_GEN
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_00 : std_logic_vector(19 downto 0) := x"029e0";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_01 : std_logic_vector(19 downto 0) := x"029f0";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_02 : std_logic_vector(19 downto 0) := x"02a00";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_03 : std_logic_vector(19 downto 0) := x"02a10";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_04 : std_logic_vector(19 downto 0) := x"02a20";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_05 : std_logic_vector(19 downto 0) := x"02a30";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_06 : std_logic_vector(19 downto 0) := x"02a40";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_07 : std_logic_vector(19 downto 0) := x"02a50";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_08 : std_logic_vector(19 downto 0) := x"02a60";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_09 : std_logic_vector(19 downto 0) := x"02a70";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_10 : std_logic_vector(19 downto 0) := x"02a80";
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_11 : std_logic_vector(19 downto 0) := x"02a90";

  --** SUPER_CHUNK_FACTOR_GEN
  constant REG_SUPER_CHUNK_FACTOR_LINK_00     : std_logic_vector(19 downto 0) := x"02de0";
  constant REG_SUPER_CHUNK_FACTOR_LINK_01     : std_logic_vector(19 downto 0) := x"02df0";
  constant REG_SUPER_CHUNK_FACTOR_LINK_02     : std_logic_vector(19 downto 0) := x"02e00";
  constant REG_SUPER_CHUNK_FACTOR_LINK_03     : std_logic_vector(19 downto 0) := x"02e10";
  constant REG_SUPER_CHUNK_FACTOR_LINK_04     : std_logic_vector(19 downto 0) := x"02e20";
  constant REG_SUPER_CHUNK_FACTOR_LINK_05     : std_logic_vector(19 downto 0) := x"02e30";
  constant REG_SUPER_CHUNK_FACTOR_LINK_06     : std_logic_vector(19 downto 0) := x"02e40";
  constant REG_SUPER_CHUNK_FACTOR_LINK_07     : std_logic_vector(19 downto 0) := x"02e50";
  constant REG_SUPER_CHUNK_FACTOR_LINK_08     : std_logic_vector(19 downto 0) := x"02e60";
  constant REG_SUPER_CHUNK_FACTOR_LINK_09     : std_logic_vector(19 downto 0) := x"02e70";
  constant REG_SUPER_CHUNK_FACTOR_LINK_10     : std_logic_vector(19 downto 0) := x"02e80";
  constant REG_SUPER_CHUNK_FACTOR_LINK_11     : std_logic_vector(19 downto 0) := x"02e90";

  --** DECODING_LINK_CB_GEN
  constant REG_DECODING_LINK_00_CB            : std_logic_vector(19 downto 0) := x"02ea0";
  constant REG_DECODING_LINK_01_CB            : std_logic_vector(19 downto 0) := x"02eb0";
  constant REG_DECODING_LINK_02_CB            : std_logic_vector(19 downto 0) := x"02ec0";
  constant REG_DECODING_LINK_03_CB            : std_logic_vector(19 downto 0) := x"02ed0";
  constant REG_DECODING_LINK_04_CB            : std_logic_vector(19 downto 0) := x"02ee0";
  constant REG_DECODING_LINK_05_CB            : std_logic_vector(19 downto 0) := x"02ef0";
  constant REG_DECODING_LINK_06_CB            : std_logic_vector(19 downto 0) := x"02f00";
  constant REG_DECODING_LINK_07_CB            : std_logic_vector(19 downto 0) := x"02f10";
  constant REG_DECODING_LINK_08_CB            : std_logic_vector(19 downto 0) := x"02f20";
  constant REG_DECODING_LINK_09_CB            : std_logic_vector(19 downto 0) := x"02f30";
  constant REG_DECODING_LINK_10_CB            : std_logic_vector(19 downto 0) := x"02f40";
  constant REG_DECODING_LINK_11_CB            : std_logic_vector(19 downto 0) := x"02f50";
  constant REG_DECODING_MASK64B66BKBLOCK      : std_logic_vector(19 downto 0) := x"02f60";
  constant REG_DECODING_DISEGROUP             : std_logic_vector(19 downto 0) := x"02f70";
  constant REG_FULLMODE_32B_SOP               : std_logic_vector(19 downto 0) := x"02f80";

  --** EncodingControlsAndMonitors
  constant REG_ENCODING_REVERSE_10B           : std_logic_vector(19 downto 0) := x"03000";

  --** ENCODING_EGROUP_CTRL_GEN

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK00_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"03010";
  constant REG_ENCODING_LINK00_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"03020";
  constant REG_ENCODING_LINK00_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"03030";
  constant REG_ENCODING_LINK00_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"03040";
  constant REG_ENCODING_LINK00_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"03050";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK01_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"03060";
  constant REG_ENCODING_LINK01_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"03070";
  constant REG_ENCODING_LINK01_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"03080";
  constant REG_ENCODING_LINK01_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"03090";
  constant REG_ENCODING_LINK01_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"030a0";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK02_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"030b0";
  constant REG_ENCODING_LINK02_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"030c0";
  constant REG_ENCODING_LINK02_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"030d0";
  constant REG_ENCODING_LINK02_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"030e0";
  constant REG_ENCODING_LINK02_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"030f0";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK03_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"03100";
  constant REG_ENCODING_LINK03_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"03110";
  constant REG_ENCODING_LINK03_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"03120";
  constant REG_ENCODING_LINK03_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"03130";
  constant REG_ENCODING_LINK03_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"03140";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK04_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"03150";
  constant REG_ENCODING_LINK04_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"03160";
  constant REG_ENCODING_LINK04_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"03170";
  constant REG_ENCODING_LINK04_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"03180";
  constant REG_ENCODING_LINK04_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"03190";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK05_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"031a0";
  constant REG_ENCODING_LINK05_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"031b0";
  constant REG_ENCODING_LINK05_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"031c0";
  constant REG_ENCODING_LINK05_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"031d0";
  constant REG_ENCODING_LINK05_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"031e0";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK06_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"031f0";
  constant REG_ENCODING_LINK06_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"03200";
  constant REG_ENCODING_LINK06_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"03210";
  constant REG_ENCODING_LINK06_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"03220";
  constant REG_ENCODING_LINK06_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"03230";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK07_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"03240";
  constant REG_ENCODING_LINK07_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"03250";
  constant REG_ENCODING_LINK07_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"03260";
  constant REG_ENCODING_LINK07_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"03270";
  constant REG_ENCODING_LINK07_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"03280";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK08_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"03290";
  constant REG_ENCODING_LINK08_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"032a0";
  constant REG_ENCODING_LINK08_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"032b0";
  constant REG_ENCODING_LINK08_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"032c0";
  constant REG_ENCODING_LINK08_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"032d0";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK09_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"032e0";
  constant REG_ENCODING_LINK09_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"032f0";
  constant REG_ENCODING_LINK09_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"03300";
  constant REG_ENCODING_LINK09_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"03310";
  constant REG_ENCODING_LINK09_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"03320";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK10_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"03330";
  constant REG_ENCODING_LINK10_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"03340";
  constant REG_ENCODING_LINK10_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"03350";
  constant REG_ENCODING_LINK10_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"03360";
  constant REG_ENCODING_LINK10_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"03370";

  --** ENCODING_EGROUP
  constant REG_ENCODING_LINK11_EGROUP0_CTRL   : std_logic_vector(19 downto 0) := x"03380";
  constant REG_ENCODING_LINK11_EGROUP1_CTRL   : std_logic_vector(19 downto 0) := x"03390";
  constant REG_ENCODING_LINK11_EGROUP2_CTRL   : std_logic_vector(19 downto 0) := x"033a0";
  constant REG_ENCODING_LINK11_EGROUP3_CTRL   : std_logic_vector(19 downto 0) := x"033b0";
  constant REG_ENCODING_LINK11_EGROUP4_CTRL   : std_logic_vector(19 downto 0) := x"033c0";

  --** MINI_EGROUP_FROMHOST_GEN
  constant REG_MINI_EGROUP_FROMHOST_00        : std_logic_vector(19 downto 0) := x"033d0";
  constant REG_MINI_EGROUP_FROMHOST_01        : std_logic_vector(19 downto 0) := x"033e0";
  constant REG_MINI_EGROUP_FROMHOST_02        : std_logic_vector(19 downto 0) := x"033f0";
  constant REG_MINI_EGROUP_FROMHOST_03        : std_logic_vector(19 downto 0) := x"03400";
  constant REG_MINI_EGROUP_FROMHOST_04        : std_logic_vector(19 downto 0) := x"03410";
  constant REG_MINI_EGROUP_FROMHOST_05        : std_logic_vector(19 downto 0) := x"03420";
  constant REG_MINI_EGROUP_FROMHOST_06        : std_logic_vector(19 downto 0) := x"03430";
  constant REG_MINI_EGROUP_FROMHOST_07        : std_logic_vector(19 downto 0) := x"03440";
  constant REG_MINI_EGROUP_FROMHOST_08        : std_logic_vector(19 downto 0) := x"03450";
  constant REG_MINI_EGROUP_FROMHOST_09        : std_logic_vector(19 downto 0) := x"03460";
  constant REG_MINI_EGROUP_FROMHOST_10        : std_logic_vector(19 downto 0) := x"03470";
  constant REG_MINI_EGROUP_FROMHOST_11        : std_logic_vector(19 downto 0) := x"03480";
  constant REG_MINI_EGROUP_FROMHOST_12        : std_logic_vector(19 downto 0) := x"03490";
  constant REG_MINI_EGROUP_FROMHOST_13        : std_logic_vector(19 downto 0) := x"034a0";
  constant REG_MINI_EGROUP_FROMHOST_14        : std_logic_vector(19 downto 0) := x"034b0";
  constant REG_MINI_EGROUP_FROMHOST_15        : std_logic_vector(19 downto 0) := x"034c0";
  constant REG_MINI_EGROUP_FROMHOST_16        : std_logic_vector(19 downto 0) := x"034d0";
  constant REG_MINI_EGROUP_FROMHOST_17        : std_logic_vector(19 downto 0) := x"034e0";
  constant REG_MINI_EGROUP_FROMHOST_18        : std_logic_vector(19 downto 0) := x"034f0";
  constant REG_MINI_EGROUP_FROMHOST_19        : std_logic_vector(19 downto 0) := x"03500";
  constant REG_MINI_EGROUP_FROMHOST_20        : std_logic_vector(19 downto 0) := x"03510";
  constant REG_MINI_EGROUP_FROMHOST_21        : std_logic_vector(19 downto 0) := x"03520";
  constant REG_MINI_EGROUP_FROMHOST_22        : std_logic_vector(19 downto 0) := x"03530";
  constant REG_MINI_EGROUP_FROMHOST_23        : std_logic_vector(19 downto 0) := x"03540";

  --** ENCODING_EGROUP_CTRL_FEI4_GEN

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03550";
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03560";
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03570";
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03580";
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03590";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"035a0";
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"035b0";
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"035c0";
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"035d0";
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"035e0";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"035f0";
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03600";
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03610";
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03620";
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03630";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03640";
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03650";
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03660";
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03670";
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03680";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03690";
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"036a0";
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"036b0";
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"036c0";
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"036d0";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"036e0";
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"036f0";
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03700";
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03710";
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03720";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03730";
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03740";
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03750";
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03760";
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03770";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03780";
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03790";
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"037a0";
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"037b0";
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"037c0";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"037d0";
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"037e0";
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"037f0";
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03800";
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03810";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03820";
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03830";
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03840";
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03850";
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03860";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03870";
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03880";
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03890";
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"038a0";
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"038b0";

  --** ENCODING_EGROUP_FEI4
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL : std_logic_vector(19 downto 0) := x"038c0";
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL : std_logic_vector(19 downto 0) := x"038d0";
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL : std_logic_vector(19 downto 0) := x"038e0";
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL : std_logic_vector(19 downto 0) := x"038f0";
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL : std_logic_vector(19 downto 0) := x"03900";

  --** YARR_DEBUG_ALLEGROUP_FROMHOST_GEN
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_00 : std_logic_vector(19 downto 0) := x"03910";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_00 : std_logic_vector(19 downto 0) := x"03920";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_01 : std_logic_vector(19 downto 0) := x"03930";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_01 : std_logic_vector(19 downto 0) := x"03940";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_02 : std_logic_vector(19 downto 0) := x"03950";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_02 : std_logic_vector(19 downto 0) := x"03960";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_03 : std_logic_vector(19 downto 0) := x"03970";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_03 : std_logic_vector(19 downto 0) := x"03980";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_04 : std_logic_vector(19 downto 0) := x"03990";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_04 : std_logic_vector(19 downto 0) := x"039a0";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_05 : std_logic_vector(19 downto 0) := x"039b0";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_05 : std_logic_vector(19 downto 0) := x"039c0";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_06 : std_logic_vector(19 downto 0) := x"039d0";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_06 : std_logic_vector(19 downto 0) := x"039e0";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_07 : std_logic_vector(19 downto 0) := x"039f0";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_07 : std_logic_vector(19 downto 0) := x"03a00";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_08 : std_logic_vector(19 downto 0) := x"03a10";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_08 : std_logic_vector(19 downto 0) := x"03a20";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_09 : std_logic_vector(19 downto 0) := x"03a30";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_09 : std_logic_vector(19 downto 0) := x"03a40";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_10 : std_logic_vector(19 downto 0) := x"03a50";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_10 : std_logic_vector(19 downto 0) := x"03a60";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_11 : std_logic_vector(19 downto 0) := x"03a70";
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_11 : std_logic_vector(19 downto 0) := x"03a80";
  constant REG_YARR_FROMHOST_CALTRIGSEQ_WE    : std_logic_vector(19 downto 0) := x"03a90";
  constant REG_YARR_FROMHOST_CALTRIGSEQ_WRDATA : std_logic_vector(19 downto 0) := x"03aa0";
  constant REG_YARR_FROMHOST_CALTRIGSEQ_WRADDR : std_logic_vector(19 downto 0) := x"03ab0";

  --** FrontendEmulatorControlsAndMonitors
  constant REG_FE_EMU_ENA                     : std_logic_vector(19 downto 0) := x"04000";
  constant REG_FE_EMU_CONFIG                  : std_logic_vector(19 downto 0) := x"04010";
  constant REG_FE_EMU_READ                    : std_logic_vector(19 downto 0) := x"04020";
  constant REG_FE_EMU_LOGIC                   : std_logic_vector(19 downto 0) := x"04030";

  --** LinkWrapperControls
  constant REG_GBT_CHANNEL_DISABLE            : std_logic_vector(19 downto 0) := x"05400";
  constant REG_GBT_GENERAL_CTRL               : std_logic_vector(19 downto 0) := x"05410";
  constant REG_GBT_MODE_CTRL                  : std_logic_vector(19 downto 0) := x"05420";
  constant REG_GBT_RXSLIDE_SELECT             : std_logic_vector(19 downto 0) := x"05480";
  constant REG_GBT_RXSLIDE_MANUAL             : std_logic_vector(19 downto 0) := x"05490";
  constant REG_GBT_TXUSRRDY                   : std_logic_vector(19 downto 0) := x"054a0";
  constant REG_GBT_RXUSRRDY                   : std_logic_vector(19 downto 0) := x"054b0";
  constant REG_GBT_SOFT_RESET                 : std_logic_vector(19 downto 0) := x"054c0";
  constant REG_GBT_GTTX_RESET                 : std_logic_vector(19 downto 0) := x"054d0";
  constant REG_GBT_GTRX_RESET                 : std_logic_vector(19 downto 0) := x"054e0";
  constant REG_GBT_PLL_RESET                  : std_logic_vector(19 downto 0) := x"054f0";
  constant REG_GBT_SOFT_TX_RESET              : std_logic_vector(19 downto 0) := x"05500";
  constant REG_GBT_SOFT_RX_RESET              : std_logic_vector(19 downto 0) := x"05510";
  constant REG_GBT_ODD_EVEN                   : std_logic_vector(19 downto 0) := x"05520";
  constant REG_GBT_TOPBOT                     : std_logic_vector(19 downto 0) := x"05530";
  constant REG_GBT_TX_TC_DLY_VALUE1           : std_logic_vector(19 downto 0) := x"05540";
  constant REG_GBT_TX_TC_DLY_VALUE2           : std_logic_vector(19 downto 0) := x"05550";
  constant REG_GBT_TX_TC_DLY_VALUE3           : std_logic_vector(19 downto 0) := x"05560";
  constant REG_GBT_TX_TC_DLY_VALUE4           : std_logic_vector(19 downto 0) := x"05570";
  constant REG_GBT_DATA_TXFORMAT1             : std_logic_vector(19 downto 0) := x"05580";
  constant REG_GBT_DATA_TXFORMAT2             : std_logic_vector(19 downto 0) := x"05590";
  constant REG_GBT_DATA_RXFORMAT1             : std_logic_vector(19 downto 0) := x"055a0";
  constant REG_GBT_DATA_RXFORMAT2             : std_logic_vector(19 downto 0) := x"055b0";
  constant REG_GBT_TX_RESET                   : std_logic_vector(19 downto 0) := x"055c0";
  constant REG_GBT_RX_RESET                   : std_logic_vector(19 downto 0) := x"055d0";
  constant REG_GBT_TX_TC_METHOD               : std_logic_vector(19 downto 0) := x"055e0";
  constant REG_GBT_OUTMUX_SEL                 : std_logic_vector(19 downto 0) := x"055f0";
  constant REG_GBT_TC_EDGE                    : std_logic_vector(19 downto 0) := x"05600";
  constant REG_GBT_TXPOLARITY                 : std_logic_vector(19 downto 0) := x"05610";
  constant REG_GBT_RXPOLARITY                 : std_logic_vector(19 downto 0) := x"05620";
  constant REG_GTH_LOOPBACK_CONTROL           : std_logic_vector(19 downto 0) := x"05630";
  constant REG_LPGBT_FEC                      : std_logic_vector(19 downto 0) := x"05640";
  constant REG_LPGBT_DATARATE                 : std_logic_vector(19 downto 0) := x"05650";
  constant REG_GBT_TOHOST_FANOUT              : std_logic_vector(19 downto 0) := x"05700";
  constant REG_GBT_TOFRONTEND_FANOUT          : std_logic_vector(19 downto 0) := x"05710";
  constant REG_FULLMODE_AUTO_RX_RESET         : std_logic_vector(19 downto 0) := x"05720";

  --** LinkWrapperMonitors
  constant REG_GBT_VERSION                    : std_logic_vector(19 downto 0) := x"06600";
  constant REG_GBT_TXRESET_DONE               : std_logic_vector(19 downto 0) := x"06680";
  constant REG_GBT_RXRESET_DONE               : std_logic_vector(19 downto 0) := x"06690";
  constant REG_GBT_TXFSMRESET_DONE            : std_logic_vector(19 downto 0) := x"066a0";
  constant REG_GBT_RXFSMRESET_DONE            : std_logic_vector(19 downto 0) := x"066b0";
  constant REG_GBT_CPLL_FBCLK_LOST            : std_logic_vector(19 downto 0) := x"066c0";
  constant REG_GBT_PLL_LOCK                   : std_logic_vector(19 downto 0) := x"066d0";
  constant REG_GBT_RXCDR_LOCK                 : std_logic_vector(19 downto 0) := x"066e0";
  constant REG_GBT_CLK_SAMPLED                : std_logic_vector(19 downto 0) := x"066f0";
  constant REG_GBT_RX_IS_HEADER               : std_logic_vector(19 downto 0) := x"06700";
  constant REG_GBT_RX_IS_DATA                 : std_logic_vector(19 downto 0) := x"06710";
  constant REG_GBT_RX_HEADER_FOUND            : std_logic_vector(19 downto 0) := x"06720";
  constant REG_GBT_ALIGNMENT_DONE             : std_logic_vector(19 downto 0) := x"06730";
  constant REG_GBT_OUT_MUX_STATUS             : std_logic_vector(19 downto 0) := x"06740";
  constant REG_GBT_ERROR                      : std_logic_vector(19 downto 0) := x"06750";
  constant REG_GBT_GBT_TOPBOT_C               : std_logic_vector(19 downto 0) := x"06760";
  constant REG_GBT_FM_RX_DISP_ERROR1          : std_logic_vector(19 downto 0) := x"06800";
  constant REG_GBT_FM_RX_DISP_ERROR2          : std_logic_vector(19 downto 0) := x"06810";
  constant REG_GBT_FM_RX_NOTINTABLE1          : std_logic_vector(19 downto 0) := x"06820";
  constant REG_GBT_FM_RX_NOTINTABLE2          : std_logic_vector(19 downto 0) := x"06830";

  --** TTCBUSYControlsAndMonitors

  --** TTC_DEC_CTRLMON
  constant REG_TTC_DEC_CTRL                   : std_logic_vector(19 downto 0) := x"07000";
  constant REG_TTC_DEC_MON                    : std_logic_vector(19 downto 0) := x"07010";

  --** TTC_BUSY_ACCEPTED_G
  constant REG_TTC_BUSY_ACCEPTED00            : std_logic_vector(19 downto 0) := x"07020";
  constant REG_TTC_BUSY_ACCEPTED01            : std_logic_vector(19 downto 0) := x"07030";
  constant REG_TTC_BUSY_ACCEPTED02            : std_logic_vector(19 downto 0) := x"07040";
  constant REG_TTC_BUSY_ACCEPTED03            : std_logic_vector(19 downto 0) := x"07050";
  constant REG_TTC_BUSY_ACCEPTED04            : std_logic_vector(19 downto 0) := x"07060";
  constant REG_TTC_BUSY_ACCEPTED05            : std_logic_vector(19 downto 0) := x"07070";
  constant REG_TTC_BUSY_ACCEPTED06            : std_logic_vector(19 downto 0) := x"07080";
  constant REG_TTC_BUSY_ACCEPTED07            : std_logic_vector(19 downto 0) := x"07090";
  constant REG_TTC_BUSY_ACCEPTED08            : std_logic_vector(19 downto 0) := x"070a0";
  constant REG_TTC_BUSY_ACCEPTED09            : std_logic_vector(19 downto 0) := x"070b0";
  constant REG_TTC_BUSY_ACCEPTED10            : std_logic_vector(19 downto 0) := x"070c0";
  constant REG_TTC_BUSY_ACCEPTED11            : std_logic_vector(19 downto 0) := x"070d0";
  constant REG_TTC_BUSY_ACCEPTED12            : std_logic_vector(19 downto 0) := x"070e0";
  constant REG_TTC_BUSY_ACCEPTED13            : std_logic_vector(19 downto 0) := x"070f0";
  constant REG_TTC_BUSY_ACCEPTED14            : std_logic_vector(19 downto 0) := x"07100";
  constant REG_TTC_BUSY_ACCEPTED15            : std_logic_vector(19 downto 0) := x"07110";
  constant REG_TTC_BUSY_ACCEPTED16            : std_logic_vector(19 downto 0) := x"07120";
  constant REG_TTC_BUSY_ACCEPTED17            : std_logic_vector(19 downto 0) := x"07130";
  constant REG_TTC_BUSY_ACCEPTED18            : std_logic_vector(19 downto 0) := x"07140";
  constant REG_TTC_BUSY_ACCEPTED19            : std_logic_vector(19 downto 0) := x"07150";
  constant REG_TTC_BUSY_ACCEPTED20            : std_logic_vector(19 downto 0) := x"07160";
  constant REG_TTC_BUSY_ACCEPTED21            : std_logic_vector(19 downto 0) := x"07170";
  constant REG_TTC_BUSY_ACCEPTED22            : std_logic_vector(19 downto 0) := x"07180";
  constant REG_TTC_BUSY_ACCEPTED23            : std_logic_vector(19 downto 0) := x"07190";
  constant REG_TTC_EMU                        : std_logic_vector(19 downto 0) := x"071a0";
  constant REG_TTC_DELAY                      : std_logic_vector(19 downto 0) := x"071b0";
  constant REG_TTC_BUSY_TIMING_CTRL           : std_logic_vector(19 downto 0) := x"074b0";
  constant REG_TTC_BUSY_CLEAR                 : std_logic_vector(19 downto 0) := x"074c0";
  constant REG_TTC_EMU_CONTROL                : std_logic_vector(19 downto 0) := x"074d0";
  constant REG_TTC_EMU_L1A_PERIOD             : std_logic_vector(19 downto 0) := x"074e0";
  constant REG_TTC_EMU_ECR_PERIOD             : std_logic_vector(19 downto 0) := x"074f0";
  constant REG_TTC_EMU_BCR_PERIOD             : std_logic_vector(19 downto 0) := x"07500";
  constant REG_TTC_EMU_LONG_CHANNEL_DATA      : std_logic_vector(19 downto 0) := x"07510";
  constant REG_TTC_EMU_RESET                  : std_logic_vector(19 downto 0) := x"07520";
  constant REG_TTC_L1ID_MONITOR               : std_logic_vector(19 downto 0) := x"07530";
  constant REG_TTC_ECR_MONITOR                : std_logic_vector(19 downto 0) := x"07540";
  constant REG_TTC_TTYPE_MONITOR              : std_logic_vector(19 downto 0) := x"07550";
  constant REG_TTC_BCR_PERIODICITY_MONITOR    : std_logic_vector(19 downto 0) := x"07560";
  constant REG_TTC_BCR_COUNTER                : std_logic_vector(19 downto 0) := x"07570";

  --** XOFF_BUSYControlsAndMonitors
  constant REG_XOFF_FM_CH_FIFO_THRESH_LOW     : std_logic_vector(19 downto 0) := x"08000";
  constant REG_XOFF_FM_CH_FIFO_THRESH_HIGH    : std_logic_vector(19 downto 0) := x"08010";
  constant REG_XOFF_FM_LOW_THRESH_CROSSED     : std_logic_vector(19 downto 0) := x"08020";
  constant REG_XOFF_FM_HIGH_THRESH            : std_logic_vector(19 downto 0) := x"08030";
  constant REG_XOFF_FM_SOFT_XOFF              : std_logic_vector(19 downto 0) := x"08040";
  constant REG_XOFF_ENABLE                    : std_logic_vector(19 downto 0) := x"08050";
  constant REG_DMA_BUSY_STATUS                : std_logic_vector(19 downto 0) := x"08060";
  constant REG_FM_BUSY_CHANNEL_STATUS         : std_logic_vector(19 downto 0) := x"08070";
  constant REG_BUSY_MAIN_OUTPUT_FIFO_THRESH   : std_logic_vector(19 downto 0) := x"08080";
  constant REG_BUSY_MAIN_OUTPUT_FIFO_STATUS   : std_logic_vector(19 downto 0) := x"08090";

  --** ELINK_BUSY_ENABLE
  constant REG_ELINK_BUSY_ENABLE00            : std_logic_vector(19 downto 0) := x"080a0";
  constant REG_ELINK_BUSY_ENABLE01            : std_logic_vector(19 downto 0) := x"080b0";
  constant REG_ELINK_BUSY_ENABLE02            : std_logic_vector(19 downto 0) := x"080c0";
  constant REG_ELINK_BUSY_ENABLE03            : std_logic_vector(19 downto 0) := x"080d0";
  constant REG_ELINK_BUSY_ENABLE04            : std_logic_vector(19 downto 0) := x"080e0";
  constant REG_ELINK_BUSY_ENABLE05            : std_logic_vector(19 downto 0) := x"080f0";
  constant REG_ELINK_BUSY_ENABLE06            : std_logic_vector(19 downto 0) := x"08100";
  constant REG_ELINK_BUSY_ENABLE07            : std_logic_vector(19 downto 0) := x"08110";
  constant REG_ELINK_BUSY_ENABLE08            : std_logic_vector(19 downto 0) := x"08120";
  constant REG_ELINK_BUSY_ENABLE09            : std_logic_vector(19 downto 0) := x"08130";
  constant REG_ELINK_BUSY_ENABLE10            : std_logic_vector(19 downto 0) := x"08140";
  constant REG_ELINK_BUSY_ENABLE11            : std_logic_vector(19 downto 0) := x"08150";
  constant REG_ELINK_BUSY_ENABLE12            : std_logic_vector(19 downto 0) := x"08160";
  constant REG_ELINK_BUSY_ENABLE13            : std_logic_vector(19 downto 0) := x"08170";
  constant REG_ELINK_BUSY_ENABLE14            : std_logic_vector(19 downto 0) := x"08180";
  constant REG_ELINK_BUSY_ENABLE15            : std_logic_vector(19 downto 0) := x"08190";
  constant REG_ELINK_BUSY_ENABLE16            : std_logic_vector(19 downto 0) := x"081a0";
  constant REG_ELINK_BUSY_ENABLE17            : std_logic_vector(19 downto 0) := x"081b0";
  constant REG_ELINK_BUSY_ENABLE18            : std_logic_vector(19 downto 0) := x"081c0";
  constant REG_ELINK_BUSY_ENABLE19            : std_logic_vector(19 downto 0) := x"081d0";
  constant REG_ELINK_BUSY_ENABLE20            : std_logic_vector(19 downto 0) := x"081e0";
  constant REG_ELINK_BUSY_ENABLE21            : std_logic_vector(19 downto 0) := x"081f0";
  constant REG_ELINK_BUSY_ENABLE22            : std_logic_vector(19 downto 0) := x"08200";
  constant REG_ELINK_BUSY_ENABLE23            : std_logic_vector(19 downto 0) := x"08210";

  --** XOFF_STATISTICS
  constant REG_XOFF_PEAK_DURATION00           : std_logic_vector(19 downto 0) := x"08220";
  constant REG_XOFF_TOTAL_DURATION00          : std_logic_vector(19 downto 0) := x"08230";
  constant REG_XOFF_COUNT00                   : std_logic_vector(19 downto 0) := x"08240";
  constant REG_XOFF_PEAK_DURATION01           : std_logic_vector(19 downto 0) := x"08250";
  constant REG_XOFF_TOTAL_DURATION01          : std_logic_vector(19 downto 0) := x"08260";
  constant REG_XOFF_COUNT01                   : std_logic_vector(19 downto 0) := x"08270";
  constant REG_XOFF_PEAK_DURATION02           : std_logic_vector(19 downto 0) := x"08280";
  constant REG_XOFF_TOTAL_DURATION02          : std_logic_vector(19 downto 0) := x"08290";
  constant REG_XOFF_COUNT02                   : std_logic_vector(19 downto 0) := x"082a0";
  constant REG_XOFF_PEAK_DURATION03           : std_logic_vector(19 downto 0) := x"082b0";
  constant REG_XOFF_TOTAL_DURATION03          : std_logic_vector(19 downto 0) := x"082c0";
  constant REG_XOFF_COUNT03                   : std_logic_vector(19 downto 0) := x"082d0";
  constant REG_XOFF_PEAK_DURATION04           : std_logic_vector(19 downto 0) := x"082e0";
  constant REG_XOFF_TOTAL_DURATION04          : std_logic_vector(19 downto 0) := x"082f0";
  constant REG_XOFF_COUNT04                   : std_logic_vector(19 downto 0) := x"08300";
  constant REG_XOFF_PEAK_DURATION05           : std_logic_vector(19 downto 0) := x"08310";
  constant REG_XOFF_TOTAL_DURATION05          : std_logic_vector(19 downto 0) := x"08320";
  constant REG_XOFF_COUNT05                   : std_logic_vector(19 downto 0) := x"08330";
  constant REG_XOFF_PEAK_DURATION06           : std_logic_vector(19 downto 0) := x"08340";
  constant REG_XOFF_TOTAL_DURATION06          : std_logic_vector(19 downto 0) := x"08350";
  constant REG_XOFF_COUNT06                   : std_logic_vector(19 downto 0) := x"08360";
  constant REG_XOFF_PEAK_DURATION07           : std_logic_vector(19 downto 0) := x"08370";
  constant REG_XOFF_TOTAL_DURATION07          : std_logic_vector(19 downto 0) := x"08380";
  constant REG_XOFF_COUNT07                   : std_logic_vector(19 downto 0) := x"08390";
  constant REG_XOFF_PEAK_DURATION08           : std_logic_vector(19 downto 0) := x"083a0";
  constant REG_XOFF_TOTAL_DURATION08          : std_logic_vector(19 downto 0) := x"083b0";
  constant REG_XOFF_COUNT08                   : std_logic_vector(19 downto 0) := x"083c0";
  constant REG_XOFF_PEAK_DURATION09           : std_logic_vector(19 downto 0) := x"083d0";
  constant REG_XOFF_TOTAL_DURATION09          : std_logic_vector(19 downto 0) := x"083e0";
  constant REG_XOFF_COUNT09                   : std_logic_vector(19 downto 0) := x"083f0";
  constant REG_XOFF_PEAK_DURATION10           : std_logic_vector(19 downto 0) := x"08400";
  constant REG_XOFF_TOTAL_DURATION10          : std_logic_vector(19 downto 0) := x"08410";
  constant REG_XOFF_COUNT10                   : std_logic_vector(19 downto 0) := x"08420";
  constant REG_XOFF_PEAK_DURATION11           : std_logic_vector(19 downto 0) := x"08430";
  constant REG_XOFF_TOTAL_DURATION11          : std_logic_vector(19 downto 0) := x"08440";
  constant REG_XOFF_COUNT11                   : std_logic_vector(19 downto 0) := x"08450";
  constant REG_XOFF_PEAK_DURATION12           : std_logic_vector(19 downto 0) := x"08460";
  constant REG_XOFF_TOTAL_DURATION12          : std_logic_vector(19 downto 0) := x"08470";
  constant REG_XOFF_COUNT12                   : std_logic_vector(19 downto 0) := x"08480";
  constant REG_XOFF_PEAK_DURATION13           : std_logic_vector(19 downto 0) := x"08490";
  constant REG_XOFF_TOTAL_DURATION13          : std_logic_vector(19 downto 0) := x"084a0";
  constant REG_XOFF_COUNT13                   : std_logic_vector(19 downto 0) := x"084b0";
  constant REG_XOFF_PEAK_DURATION14           : std_logic_vector(19 downto 0) := x"084c0";
  constant REG_XOFF_TOTAL_DURATION14          : std_logic_vector(19 downto 0) := x"084d0";
  constant REG_XOFF_COUNT14                   : std_logic_vector(19 downto 0) := x"084e0";
  constant REG_XOFF_PEAK_DURATION15           : std_logic_vector(19 downto 0) := x"084f0";
  constant REG_XOFF_TOTAL_DURATION15          : std_logic_vector(19 downto 0) := x"08500";
  constant REG_XOFF_COUNT15                   : std_logic_vector(19 downto 0) := x"08510";
  constant REG_XOFF_PEAK_DURATION16           : std_logic_vector(19 downto 0) := x"08520";
  constant REG_XOFF_TOTAL_DURATION16          : std_logic_vector(19 downto 0) := x"08530";
  constant REG_XOFF_COUNT16                   : std_logic_vector(19 downto 0) := x"08540";
  constant REG_XOFF_PEAK_DURATION17           : std_logic_vector(19 downto 0) := x"08550";
  constant REG_XOFF_TOTAL_DURATION17          : std_logic_vector(19 downto 0) := x"08560";
  constant REG_XOFF_COUNT17                   : std_logic_vector(19 downto 0) := x"08570";
  constant REG_XOFF_PEAK_DURATION18           : std_logic_vector(19 downto 0) := x"08580";
  constant REG_XOFF_TOTAL_DURATION18          : std_logic_vector(19 downto 0) := x"08590";
  constant REG_XOFF_COUNT18                   : std_logic_vector(19 downto 0) := x"085a0";
  constant REG_XOFF_PEAK_DURATION19           : std_logic_vector(19 downto 0) := x"085b0";
  constant REG_XOFF_TOTAL_DURATION19          : std_logic_vector(19 downto 0) := x"085c0";
  constant REG_XOFF_COUNT19                   : std_logic_vector(19 downto 0) := x"085d0";
  constant REG_XOFF_PEAK_DURATION20           : std_logic_vector(19 downto 0) := x"085e0";
  constant REG_XOFF_TOTAL_DURATION20          : std_logic_vector(19 downto 0) := x"085f0";
  constant REG_XOFF_COUNT20                   : std_logic_vector(19 downto 0) := x"08600";
  constant REG_XOFF_PEAK_DURATION21           : std_logic_vector(19 downto 0) := x"08610";
  constant REG_XOFF_TOTAL_DURATION21          : std_logic_vector(19 downto 0) := x"08620";
  constant REG_XOFF_COUNT21                   : std_logic_vector(19 downto 0) := x"08630";
  constant REG_XOFF_PEAK_DURATION22           : std_logic_vector(19 downto 0) := x"08640";
  constant REG_XOFF_TOTAL_DURATION22          : std_logic_vector(19 downto 0) := x"08650";
  constant REG_XOFF_COUNT22                   : std_logic_vector(19 downto 0) := x"08660";
  constant REG_XOFF_PEAK_DURATION23           : std_logic_vector(19 downto 0) := x"08670";
  constant REG_XOFF_TOTAL_DURATION23          : std_logic_vector(19 downto 0) := x"08680";
  constant REG_XOFF_COUNT23                   : std_logic_vector(19 downto 0) := x"08690";
  constant REG_BUSY_TOHOST_ENABLE             : std_logic_vector(19 downto 0) := x"086a0";

  --** HouseKeepingControlsAndMonitors
  constant REG_HK_CTRL_I2C                    : std_logic_vector(19 downto 0) := x"09000";
  constant REG_HK_CTRL_FMC                    : std_logic_vector(19 downto 0) := x"09010";
  constant REG_HK_MON_FMC                     : std_logic_vector(19 downto 0) := x"09020";
  constant REG_MMCM_MAIN                      : std_logic_vector(19 downto 0) := x"09300";
  constant REG_LMK_LOCKED                     : std_logic_vector(19 downto 0) := x"09310";
  constant REG_FPGA_CORE_TEMP                 : std_logic_vector(19 downto 0) := x"09320";
  constant REG_FPGA_CORE_VCCINT               : std_logic_vector(19 downto 0) := x"09330";
  constant REG_FPGA_CORE_VCCAUX               : std_logic_vector(19 downto 0) := x"09340";
  constant REG_FPGA_CORE_VCCBRAM              : std_logic_vector(19 downto 0) := x"09350";
  constant REG_FPGA_DNA                       : std_logic_vector(19 downto 0) := x"09360";
  constant REG_I2C_WR                         : std_logic_vector(19 downto 0) := x"09420";
  constant REG_I2C_RD                         : std_logic_vector(19 downto 0) := x"09430";
  constant REG_INT_TEST                       : std_logic_vector(19 downto 0) := x"09800";
  constant REG_CONFIG_FLASH_WR                : std_logic_vector(19 downto 0) := x"09810";
  constant REG_CONFIG_FLASH_RD                : std_logic_vector(19 downto 0) := x"09820";
  constant REG_SI5324_STATUS                  : std_logic_vector(19 downto 0) := x"09830";
  constant REG_TACH_CNT                       : std_logic_vector(19 downto 0) := x"09840";
  constant REG_RXUSRCLK_FREQ                  : std_logic_vector(19 downto 0) := x"09850";

  --** Generators
  constant REG_FELIG_L1ID_RESET               : std_logic_vector(19 downto 0) := x"0a000";

  --** FELIG_DATA_GEN_CONFIG_ARR
  constant REG_FELIG_DATA_GEN_CONFIG_00       : std_logic_vector(19 downto 0) := x"0a020";
  constant REG_FELIG_DATA_GEN_CONFIG_01       : std_logic_vector(19 downto 0) := x"0a030";
  constant REG_FELIG_DATA_GEN_CONFIG_02       : std_logic_vector(19 downto 0) := x"0a040";
  constant REG_FELIG_DATA_GEN_CONFIG_03       : std_logic_vector(19 downto 0) := x"0a050";
  constant REG_FELIG_DATA_GEN_CONFIG_04       : std_logic_vector(19 downto 0) := x"0a060";
  constant REG_FELIG_DATA_GEN_CONFIG_05       : std_logic_vector(19 downto 0) := x"0a070";
  constant REG_FELIG_DATA_GEN_CONFIG_06       : std_logic_vector(19 downto 0) := x"0a080";
  constant REG_FELIG_DATA_GEN_CONFIG_07       : std_logic_vector(19 downto 0) := x"0a090";
  constant REG_FELIG_DATA_GEN_CONFIG_08       : std_logic_vector(19 downto 0) := x"0a0a0";
  constant REG_FELIG_DATA_GEN_CONFIG_09       : std_logic_vector(19 downto 0) := x"0a0b0";
  constant REG_FELIG_DATA_GEN_CONFIG_10       : std_logic_vector(19 downto 0) := x"0a0c0";
  constant REG_FELIG_DATA_GEN_CONFIG_11       : std_logic_vector(19 downto 0) := x"0a0d0";
  constant REG_FELIG_DATA_GEN_CONFIG_12       : std_logic_vector(19 downto 0) := x"0a0e0";
  constant REG_FELIG_DATA_GEN_CONFIG_13       : std_logic_vector(19 downto 0) := x"0a0f0";
  constant REG_FELIG_DATA_GEN_CONFIG_14       : std_logic_vector(19 downto 0) := x"0a100";
  constant REG_FELIG_DATA_GEN_CONFIG_15       : std_logic_vector(19 downto 0) := x"0a110";
  constant REG_FELIG_DATA_GEN_CONFIG_16       : std_logic_vector(19 downto 0) := x"0a120";
  constant REG_FELIG_DATA_GEN_CONFIG_17       : std_logic_vector(19 downto 0) := x"0a130";
  constant REG_FELIG_DATA_GEN_CONFIG_18       : std_logic_vector(19 downto 0) := x"0a140";
  constant REG_FELIG_DATA_GEN_CONFIG_19       : std_logic_vector(19 downto 0) := x"0a150";
  constant REG_FELIG_DATA_GEN_CONFIG_20       : std_logic_vector(19 downto 0) := x"0a160";
  constant REG_FELIG_DATA_GEN_CONFIG_21       : std_logic_vector(19 downto 0) := x"0a170";
  constant REG_FELIG_DATA_GEN_CONFIG_22       : std_logic_vector(19 downto 0) := x"0a180";
  constant REG_FELIG_DATA_GEN_CONFIG_23       : std_logic_vector(19 downto 0) := x"0a190";

  --** FELIG_ELINK_CONFIG_ARR
  constant REG_FELIG_ELINK_CONFIG_00          : std_logic_vector(19 downto 0) := x"0a1a0";
  constant REG_FELIG_ELINK_CONFIG_01          : std_logic_vector(19 downto 0) := x"0a1b0";
  constant REG_FELIG_ELINK_CONFIG_02          : std_logic_vector(19 downto 0) := x"0a1c0";
  constant REG_FELIG_ELINK_CONFIG_03          : std_logic_vector(19 downto 0) := x"0a1d0";
  constant REG_FELIG_ELINK_CONFIG_04          : std_logic_vector(19 downto 0) := x"0a1e0";
  constant REG_FELIG_ELINK_CONFIG_05          : std_logic_vector(19 downto 0) := x"0a1f0";
  constant REG_FELIG_ELINK_CONFIG_06          : std_logic_vector(19 downto 0) := x"0a200";
  constant REG_FELIG_ELINK_CONFIG_07          : std_logic_vector(19 downto 0) := x"0a210";
  constant REG_FELIG_ELINK_CONFIG_08          : std_logic_vector(19 downto 0) := x"0a220";
  constant REG_FELIG_ELINK_CONFIG_09          : std_logic_vector(19 downto 0) := x"0a230";
  constant REG_FELIG_ELINK_CONFIG_10          : std_logic_vector(19 downto 0) := x"0a240";
  constant REG_FELIG_ELINK_CONFIG_11          : std_logic_vector(19 downto 0) := x"0a250";
  constant REG_FELIG_ELINK_CONFIG_12          : std_logic_vector(19 downto 0) := x"0a260";
  constant REG_FELIG_ELINK_CONFIG_13          : std_logic_vector(19 downto 0) := x"0a270";
  constant REG_FELIG_ELINK_CONFIG_14          : std_logic_vector(19 downto 0) := x"0a280";
  constant REG_FELIG_ELINK_CONFIG_15          : std_logic_vector(19 downto 0) := x"0a290";
  constant REG_FELIG_ELINK_CONFIG_16          : std_logic_vector(19 downto 0) := x"0a2a0";
  constant REG_FELIG_ELINK_CONFIG_17          : std_logic_vector(19 downto 0) := x"0a2b0";
  constant REG_FELIG_ELINK_CONFIG_18          : std_logic_vector(19 downto 0) := x"0a2c0";
  constant REG_FELIG_ELINK_CONFIG_19          : std_logic_vector(19 downto 0) := x"0a2d0";
  constant REG_FELIG_ELINK_CONFIG_20          : std_logic_vector(19 downto 0) := x"0a2e0";
  constant REG_FELIG_ELINK_CONFIG_21          : std_logic_vector(19 downto 0) := x"0a2f0";
  constant REG_FELIG_ELINK_CONFIG_22          : std_logic_vector(19 downto 0) := x"0a300";
  constant REG_FELIG_ELINK_CONFIG_23          : std_logic_vector(19 downto 0) := x"0a310";

  --** FELIG_ELINK_ENABLE_ARR
  constant REG_FELIG_ELINK_ENABLE_00          : std_logic_vector(19 downto 0) := x"0a320";
  constant REG_FELIG_ELINK_ENABLE_01          : std_logic_vector(19 downto 0) := x"0a330";
  constant REG_FELIG_ELINK_ENABLE_02          : std_logic_vector(19 downto 0) := x"0a340";
  constant REG_FELIG_ELINK_ENABLE_03          : std_logic_vector(19 downto 0) := x"0a350";
  constant REG_FELIG_ELINK_ENABLE_04          : std_logic_vector(19 downto 0) := x"0a360";
  constant REG_FELIG_ELINK_ENABLE_05          : std_logic_vector(19 downto 0) := x"0a370";
  constant REG_FELIG_ELINK_ENABLE_06          : std_logic_vector(19 downto 0) := x"0a380";
  constant REG_FELIG_ELINK_ENABLE_07          : std_logic_vector(19 downto 0) := x"0a390";
  constant REG_FELIG_ELINK_ENABLE_08          : std_logic_vector(19 downto 0) := x"0a3a0";
  constant REG_FELIG_ELINK_ENABLE_09          : std_logic_vector(19 downto 0) := x"0a3b0";
  constant REG_FELIG_ELINK_ENABLE_10          : std_logic_vector(19 downto 0) := x"0a3c0";
  constant REG_FELIG_ELINK_ENABLE_11          : std_logic_vector(19 downto 0) := x"0a3d0";
  constant REG_FELIG_ELINK_ENABLE_12          : std_logic_vector(19 downto 0) := x"0a3e0";
  constant REG_FELIG_ELINK_ENABLE_13          : std_logic_vector(19 downto 0) := x"0a3f0";
  constant REG_FELIG_ELINK_ENABLE_14          : std_logic_vector(19 downto 0) := x"0a400";
  constant REG_FELIG_ELINK_ENABLE_15          : std_logic_vector(19 downto 0) := x"0a410";
  constant REG_FELIG_ELINK_ENABLE_16          : std_logic_vector(19 downto 0) := x"0a420";
  constant REG_FELIG_ELINK_ENABLE_17          : std_logic_vector(19 downto 0) := x"0a430";
  constant REG_FELIG_ELINK_ENABLE_18          : std_logic_vector(19 downto 0) := x"0a440";
  constant REG_FELIG_ELINK_ENABLE_19          : std_logic_vector(19 downto 0) := x"0a450";
  constant REG_FELIG_ELINK_ENABLE_20          : std_logic_vector(19 downto 0) := x"0a460";
  constant REG_FELIG_ELINK_ENABLE_21          : std_logic_vector(19 downto 0) := x"0a470";
  constant REG_FELIG_ELINK_ENABLE_22          : std_logic_vector(19 downto 0) := x"0a480";
  constant REG_FELIG_ELINK_ENABLE_23          : std_logic_vector(19 downto 0) := x"0a490";
  constant REG_FELIG_GLOBAL_CONTROL           : std_logic_vector(19 downto 0) := x"0a4a0";

  --** FELIG_LANE_CONFIG_ARR
  constant REG_FELIG_LANE_CONFIG_00           : std_logic_vector(19 downto 0) := x"0a4b0";
  constant REG_FELIG_LANE_CONFIG_01           : std_logic_vector(19 downto 0) := x"0a4c0";
  constant REG_FELIG_LANE_CONFIG_02           : std_logic_vector(19 downto 0) := x"0a4d0";
  constant REG_FELIG_LANE_CONFIG_03           : std_logic_vector(19 downto 0) := x"0a4e0";
  constant REG_FELIG_LANE_CONFIG_04           : std_logic_vector(19 downto 0) := x"0a4f0";
  constant REG_FELIG_LANE_CONFIG_05           : std_logic_vector(19 downto 0) := x"0a500";
  constant REG_FELIG_LANE_CONFIG_06           : std_logic_vector(19 downto 0) := x"0a510";
  constant REG_FELIG_LANE_CONFIG_07           : std_logic_vector(19 downto 0) := x"0a520";
  constant REG_FELIG_LANE_CONFIG_08           : std_logic_vector(19 downto 0) := x"0a530";
  constant REG_FELIG_LANE_CONFIG_09           : std_logic_vector(19 downto 0) := x"0a540";
  constant REG_FELIG_LANE_CONFIG_10           : std_logic_vector(19 downto 0) := x"0a550";
  constant REG_FELIG_LANE_CONFIG_11           : std_logic_vector(19 downto 0) := x"0a560";
  constant REG_FELIG_LANE_CONFIG_12           : std_logic_vector(19 downto 0) := x"0a570";
  constant REG_FELIG_LANE_CONFIG_13           : std_logic_vector(19 downto 0) := x"0a580";
  constant REG_FELIG_LANE_CONFIG_14           : std_logic_vector(19 downto 0) := x"0a590";
  constant REG_FELIG_LANE_CONFIG_15           : std_logic_vector(19 downto 0) := x"0a5a0";
  constant REG_FELIG_LANE_CONFIG_16           : std_logic_vector(19 downto 0) := x"0a5b0";
  constant REG_FELIG_LANE_CONFIG_17           : std_logic_vector(19 downto 0) := x"0a5c0";
  constant REG_FELIG_LANE_CONFIG_18           : std_logic_vector(19 downto 0) := x"0a5d0";
  constant REG_FELIG_LANE_CONFIG_19           : std_logic_vector(19 downto 0) := x"0a5e0";
  constant REG_FELIG_LANE_CONFIG_20           : std_logic_vector(19 downto 0) := x"0a5f0";
  constant REG_FELIG_LANE_CONFIG_21           : std_logic_vector(19 downto 0) := x"0a600";
  constant REG_FELIG_LANE_CONFIG_22           : std_logic_vector(19 downto 0) := x"0a610";
  constant REG_FELIG_LANE_CONFIG_23           : std_logic_vector(19 downto 0) := x"0a620";

  --** FELIG_MON_TTC_0_ARR
  constant REG_FELIG_MON_TTC_0_00             : std_logic_vector(19 downto 0) := x"0a630";
  constant REG_FELIG_MON_TTC_0_01             : std_logic_vector(19 downto 0) := x"0a640";
  constant REG_FELIG_MON_TTC_0_02             : std_logic_vector(19 downto 0) := x"0a650";
  constant REG_FELIG_MON_TTC_0_03             : std_logic_vector(19 downto 0) := x"0a660";
  constant REG_FELIG_MON_TTC_0_04             : std_logic_vector(19 downto 0) := x"0a670";
  constant REG_FELIG_MON_TTC_0_05             : std_logic_vector(19 downto 0) := x"0a680";
  constant REG_FELIG_MON_TTC_0_06             : std_logic_vector(19 downto 0) := x"0a690";
  constant REG_FELIG_MON_TTC_0_07             : std_logic_vector(19 downto 0) := x"0a6a0";
  constant REG_FELIG_MON_TTC_0_08             : std_logic_vector(19 downto 0) := x"0a6b0";
  constant REG_FELIG_MON_TTC_0_09             : std_logic_vector(19 downto 0) := x"0a6c0";
  constant REG_FELIG_MON_TTC_0_10             : std_logic_vector(19 downto 0) := x"0a6d0";
  constant REG_FELIG_MON_TTC_0_11             : std_logic_vector(19 downto 0) := x"0a6e0";
  constant REG_FELIG_MON_TTC_0_12             : std_logic_vector(19 downto 0) := x"0a6f0";
  constant REG_FELIG_MON_TTC_0_13             : std_logic_vector(19 downto 0) := x"0a700";
  constant REG_FELIG_MON_TTC_0_14             : std_logic_vector(19 downto 0) := x"0a710";
  constant REG_FELIG_MON_TTC_0_15             : std_logic_vector(19 downto 0) := x"0a720";
  constant REG_FELIG_MON_TTC_0_16             : std_logic_vector(19 downto 0) := x"0a730";
  constant REG_FELIG_MON_TTC_0_17             : std_logic_vector(19 downto 0) := x"0a740";
  constant REG_FELIG_MON_TTC_0_18             : std_logic_vector(19 downto 0) := x"0a750";
  constant REG_FELIG_MON_TTC_0_19             : std_logic_vector(19 downto 0) := x"0a760";
  constant REG_FELIG_MON_TTC_0_20             : std_logic_vector(19 downto 0) := x"0a770";
  constant REG_FELIG_MON_TTC_0_21             : std_logic_vector(19 downto 0) := x"0a780";
  constant REG_FELIG_MON_TTC_0_22             : std_logic_vector(19 downto 0) := x"0a790";
  constant REG_FELIG_MON_TTC_0_23             : std_logic_vector(19 downto 0) := x"0a7a0";

  --** FELIG_MON_TTC_1_ARR
  constant REG_FELIG_MON_TTC_1_00             : std_logic_vector(19 downto 0) := x"0a7b0";
  constant REG_FELIG_MON_TTC_1_01             : std_logic_vector(19 downto 0) := x"0a7c0";
  constant REG_FELIG_MON_TTC_1_02             : std_logic_vector(19 downto 0) := x"0a7d0";
  constant REG_FELIG_MON_TTC_1_03             : std_logic_vector(19 downto 0) := x"0a7e0";
  constant REG_FELIG_MON_TTC_1_04             : std_logic_vector(19 downto 0) := x"0a7f0";
  constant REG_FELIG_MON_TTC_1_05             : std_logic_vector(19 downto 0) := x"0a800";
  constant REG_FELIG_MON_TTC_1_06             : std_logic_vector(19 downto 0) := x"0a810";
  constant REG_FELIG_MON_TTC_1_07             : std_logic_vector(19 downto 0) := x"0a820";
  constant REG_FELIG_MON_TTC_1_08             : std_logic_vector(19 downto 0) := x"0a830";
  constant REG_FELIG_MON_TTC_1_09             : std_logic_vector(19 downto 0) := x"0a840";
  constant REG_FELIG_MON_TTC_1_10             : std_logic_vector(19 downto 0) := x"0a850";
  constant REG_FELIG_MON_TTC_1_11             : std_logic_vector(19 downto 0) := x"0a860";
  constant REG_FELIG_MON_TTC_1_12             : std_logic_vector(19 downto 0) := x"0a870";
  constant REG_FELIG_MON_TTC_1_13             : std_logic_vector(19 downto 0) := x"0a880";
  constant REG_FELIG_MON_TTC_1_14             : std_logic_vector(19 downto 0) := x"0a890";
  constant REG_FELIG_MON_TTC_1_15             : std_logic_vector(19 downto 0) := x"0a8a0";
  constant REG_FELIG_MON_TTC_1_16             : std_logic_vector(19 downto 0) := x"0a8b0";
  constant REG_FELIG_MON_TTC_1_17             : std_logic_vector(19 downto 0) := x"0a8c0";
  constant REG_FELIG_MON_TTC_1_18             : std_logic_vector(19 downto 0) := x"0a8d0";
  constant REG_FELIG_MON_TTC_1_19             : std_logic_vector(19 downto 0) := x"0a8e0";
  constant REG_FELIG_MON_TTC_1_20             : std_logic_vector(19 downto 0) := x"0a8f0";
  constant REG_FELIG_MON_TTC_1_21             : std_logic_vector(19 downto 0) := x"0a900";
  constant REG_FELIG_MON_TTC_1_22             : std_logic_vector(19 downto 0) := x"0a910";
  constant REG_FELIG_MON_TTC_1_23             : std_logic_vector(19 downto 0) := x"0a920";

  --** FELIG_MON_COUNTERS_ARR
  constant REG_FELIG_MON_COUNTERS_00          : std_logic_vector(19 downto 0) := x"0a930";
  constant REG_FELIG_MON_COUNTERS_01          : std_logic_vector(19 downto 0) := x"0a940";
  constant REG_FELIG_MON_COUNTERS_02          : std_logic_vector(19 downto 0) := x"0a950";
  constant REG_FELIG_MON_COUNTERS_03          : std_logic_vector(19 downto 0) := x"0a960";
  constant REG_FELIG_MON_COUNTERS_04          : std_logic_vector(19 downto 0) := x"0a970";
  constant REG_FELIG_MON_COUNTERS_05          : std_logic_vector(19 downto 0) := x"0a980";
  constant REG_FELIG_MON_COUNTERS_06          : std_logic_vector(19 downto 0) := x"0a990";
  constant REG_FELIG_MON_COUNTERS_07          : std_logic_vector(19 downto 0) := x"0a9a0";
  constant REG_FELIG_MON_COUNTERS_08          : std_logic_vector(19 downto 0) := x"0a9b0";
  constant REG_FELIG_MON_COUNTERS_09          : std_logic_vector(19 downto 0) := x"0a9c0";
  constant REG_FELIG_MON_COUNTERS_10          : std_logic_vector(19 downto 0) := x"0a9d0";
  constant REG_FELIG_MON_COUNTERS_11          : std_logic_vector(19 downto 0) := x"0a9e0";
  constant REG_FELIG_MON_COUNTERS_12          : std_logic_vector(19 downto 0) := x"0a9f0";
  constant REG_FELIG_MON_COUNTERS_13          : std_logic_vector(19 downto 0) := x"0aa00";
  constant REG_FELIG_MON_COUNTERS_14          : std_logic_vector(19 downto 0) := x"0aa10";
  constant REG_FELIG_MON_COUNTERS_15          : std_logic_vector(19 downto 0) := x"0aa20";
  constant REG_FELIG_MON_COUNTERS_16          : std_logic_vector(19 downto 0) := x"0aa30";
  constant REG_FELIG_MON_COUNTERS_17          : std_logic_vector(19 downto 0) := x"0aa40";
  constant REG_FELIG_MON_COUNTERS_18          : std_logic_vector(19 downto 0) := x"0aa50";
  constant REG_FELIG_MON_COUNTERS_19          : std_logic_vector(19 downto 0) := x"0aa60";
  constant REG_FELIG_MON_COUNTERS_20          : std_logic_vector(19 downto 0) := x"0aa70";
  constant REG_FELIG_MON_COUNTERS_21          : std_logic_vector(19 downto 0) := x"0aa80";
  constant REG_FELIG_MON_COUNTERS_22          : std_logic_vector(19 downto 0) := x"0aa90";
  constant REG_FELIG_MON_COUNTERS_23          : std_logic_vector(19 downto 0) := x"0aaa0";

  --** FELIG_MON_FREQ_ARR
  constant REG_FELIG_MON_FREQ_00              : std_logic_vector(19 downto 0) := x"0aab0";
  constant REG_FELIG_MON_FREQ_01              : std_logic_vector(19 downto 0) := x"0aac0";
  constant REG_FELIG_MON_FREQ_02              : std_logic_vector(19 downto 0) := x"0aad0";
  constant REG_FELIG_MON_FREQ_03              : std_logic_vector(19 downto 0) := x"0aae0";
  constant REG_FELIG_MON_FREQ_04              : std_logic_vector(19 downto 0) := x"0aaf0";
  constant REG_FELIG_MON_FREQ_05              : std_logic_vector(19 downto 0) := x"0ab00";
  constant REG_FELIG_MON_FREQ_06              : std_logic_vector(19 downto 0) := x"0ab10";
  constant REG_FELIG_MON_FREQ_07              : std_logic_vector(19 downto 0) := x"0ab20";
  constant REG_FELIG_MON_FREQ_08              : std_logic_vector(19 downto 0) := x"0ab30";
  constant REG_FELIG_MON_FREQ_09              : std_logic_vector(19 downto 0) := x"0ab40";
  constant REG_FELIG_MON_FREQ_10              : std_logic_vector(19 downto 0) := x"0ab50";
  constant REG_FELIG_MON_FREQ_11              : std_logic_vector(19 downto 0) := x"0ab60";
  constant REG_FELIG_MON_FREQ_12              : std_logic_vector(19 downto 0) := x"0ab70";
  constant REG_FELIG_MON_FREQ_13              : std_logic_vector(19 downto 0) := x"0ab80";
  constant REG_FELIG_MON_FREQ_14              : std_logic_vector(19 downto 0) := x"0ab90";
  constant REG_FELIG_MON_FREQ_15              : std_logic_vector(19 downto 0) := x"0aba0";
  constant REG_FELIG_MON_FREQ_16              : std_logic_vector(19 downto 0) := x"0abb0";
  constant REG_FELIG_MON_FREQ_17              : std_logic_vector(19 downto 0) := x"0abc0";
  constant REG_FELIG_MON_FREQ_18              : std_logic_vector(19 downto 0) := x"0abd0";
  constant REG_FELIG_MON_FREQ_19              : std_logic_vector(19 downto 0) := x"0abe0";
  constant REG_FELIG_MON_FREQ_20              : std_logic_vector(19 downto 0) := x"0abf0";
  constant REG_FELIG_MON_FREQ_21              : std_logic_vector(19 downto 0) := x"0ac00";
  constant REG_FELIG_MON_FREQ_22              : std_logic_vector(19 downto 0) := x"0ac10";
  constant REG_FELIG_MON_FREQ_23              : std_logic_vector(19 downto 0) := x"0ac20";
  constant REG_FELIG_MON_FREQ_GLOBAL          : std_logic_vector(19 downto 0) := x"0ac30";

  --** FELIG_MON_L1A_ID_ARR
  constant REG_FELIG_MON_L1A_ID_00            : std_logic_vector(19 downto 0) := x"0ac40";
  constant REG_FELIG_MON_L1A_ID_01            : std_logic_vector(19 downto 0) := x"0ac50";
  constant REG_FELIG_MON_L1A_ID_02            : std_logic_vector(19 downto 0) := x"0ac60";
  constant REG_FELIG_MON_L1A_ID_03            : std_logic_vector(19 downto 0) := x"0ac70";
  constant REG_FELIG_MON_L1A_ID_04            : std_logic_vector(19 downto 0) := x"0ac80";
  constant REG_FELIG_MON_L1A_ID_05            : std_logic_vector(19 downto 0) := x"0ac90";
  constant REG_FELIG_MON_L1A_ID_06            : std_logic_vector(19 downto 0) := x"0aca0";
  constant REG_FELIG_MON_L1A_ID_07            : std_logic_vector(19 downto 0) := x"0acb0";
  constant REG_FELIG_MON_L1A_ID_08            : std_logic_vector(19 downto 0) := x"0acc0";
  constant REG_FELIG_MON_L1A_ID_09            : std_logic_vector(19 downto 0) := x"0acd0";
  constant REG_FELIG_MON_L1A_ID_10            : std_logic_vector(19 downto 0) := x"0ace0";
  constant REG_FELIG_MON_L1A_ID_11            : std_logic_vector(19 downto 0) := x"0acf0";
  constant REG_FELIG_MON_L1A_ID_12            : std_logic_vector(19 downto 0) := x"0ad00";
  constant REG_FELIG_MON_L1A_ID_13            : std_logic_vector(19 downto 0) := x"0ad10";
  constant REG_FELIG_MON_L1A_ID_14            : std_logic_vector(19 downto 0) := x"0ad20";
  constant REG_FELIG_MON_L1A_ID_15            : std_logic_vector(19 downto 0) := x"0ad30";
  constant REG_FELIG_MON_L1A_ID_16            : std_logic_vector(19 downto 0) := x"0ad40";
  constant REG_FELIG_MON_L1A_ID_17            : std_logic_vector(19 downto 0) := x"0ad50";
  constant REG_FELIG_MON_L1A_ID_18            : std_logic_vector(19 downto 0) := x"0ad60";
  constant REG_FELIG_MON_L1A_ID_19            : std_logic_vector(19 downto 0) := x"0ad70";
  constant REG_FELIG_MON_L1A_ID_20            : std_logic_vector(19 downto 0) := x"0ad80";
  constant REG_FELIG_MON_L1A_ID_21            : std_logic_vector(19 downto 0) := x"0ad90";
  constant REG_FELIG_MON_L1A_ID_22            : std_logic_vector(19 downto 0) := x"0ada0";
  constant REG_FELIG_MON_L1A_ID_23            : std_logic_vector(19 downto 0) := x"0adb0";

  --** FELIG_MON_PICXO_ARR
  constant REG_FELIG_MON_PICXO_00             : std_logic_vector(19 downto 0) := x"0adc0";
  constant REG_FELIG_MON_PICXO_01             : std_logic_vector(19 downto 0) := x"0add0";
  constant REG_FELIG_MON_PICXO_02             : std_logic_vector(19 downto 0) := x"0ade0";
  constant REG_FELIG_MON_PICXO_03             : std_logic_vector(19 downto 0) := x"0adf0";
  constant REG_FELIG_MON_PICXO_04             : std_logic_vector(19 downto 0) := x"0ae00";
  constant REG_FELIG_MON_PICXO_05             : std_logic_vector(19 downto 0) := x"0ae10";
  constant REG_FELIG_MON_PICXO_06             : std_logic_vector(19 downto 0) := x"0ae20";
  constant REG_FELIG_MON_PICXO_07             : std_logic_vector(19 downto 0) := x"0ae30";
  constant REG_FELIG_MON_PICXO_08             : std_logic_vector(19 downto 0) := x"0ae40";
  constant REG_FELIG_MON_PICXO_09             : std_logic_vector(19 downto 0) := x"0ae50";
  constant REG_FELIG_MON_PICXO_10             : std_logic_vector(19 downto 0) := x"0ae60";
  constant REG_FELIG_MON_PICXO_11             : std_logic_vector(19 downto 0) := x"0ae70";
  constant REG_FELIG_MON_PICXO_12             : std_logic_vector(19 downto 0) := x"0ae80";
  constant REG_FELIG_MON_PICXO_13             : std_logic_vector(19 downto 0) := x"0ae90";
  constant REG_FELIG_MON_PICXO_14             : std_logic_vector(19 downto 0) := x"0aea0";
  constant REG_FELIG_MON_PICXO_15             : std_logic_vector(19 downto 0) := x"0aeb0";
  constant REG_FELIG_MON_PICXO_16             : std_logic_vector(19 downto 0) := x"0aec0";
  constant REG_FELIG_MON_PICXO_17             : std_logic_vector(19 downto 0) := x"0aed0";
  constant REG_FELIG_MON_PICXO_18             : std_logic_vector(19 downto 0) := x"0aee0";
  constant REG_FELIG_MON_PICXO_19             : std_logic_vector(19 downto 0) := x"0aef0";
  constant REG_FELIG_MON_PICXO_20             : std_logic_vector(19 downto 0) := x"0af00";
  constant REG_FELIG_MON_PICXO_21             : std_logic_vector(19 downto 0) := x"0af10";
  constant REG_FELIG_MON_PICXO_22             : std_logic_vector(19 downto 0) := x"0af20";
  constant REG_FELIG_MON_PICXO_23             : std_logic_vector(19 downto 0) := x"0af30";
  constant REG_FELIG_RESET                    : std_logic_vector(19 downto 0) := x"0af40";
  constant REG_FELIG_RX_SLIDE_RESET           : std_logic_vector(19 downto 0) := x"0af50";

  --** FELIG_ITK_STRIPS_DATA_GEN_CONFIG_ARR
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_00 : std_logic_vector(19 downto 0) := x"0af60";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_01 : std_logic_vector(19 downto 0) := x"0af70";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_02 : std_logic_vector(19 downto 0) := x"0af80";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_03 : std_logic_vector(19 downto 0) := x"0af90";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_04 : std_logic_vector(19 downto 0) := x"0afa0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_05 : std_logic_vector(19 downto 0) := x"0afb0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_06 : std_logic_vector(19 downto 0) := x"0afc0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_07 : std_logic_vector(19 downto 0) := x"0afd0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_08 : std_logic_vector(19 downto 0) := x"0afe0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_09 : std_logic_vector(19 downto 0) := x"0aff0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_10 : std_logic_vector(19 downto 0) := x"0b000";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_11 : std_logic_vector(19 downto 0) := x"0b010";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_12 : std_logic_vector(19 downto 0) := x"0b020";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_13 : std_logic_vector(19 downto 0) := x"0b030";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_14 : std_logic_vector(19 downto 0) := x"0b040";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_15 : std_logic_vector(19 downto 0) := x"0b050";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_16 : std_logic_vector(19 downto 0) := x"0b060";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_17 : std_logic_vector(19 downto 0) := x"0b070";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_18 : std_logic_vector(19 downto 0) := x"0b080";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_19 : std_logic_vector(19 downto 0) := x"0b090";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_20 : std_logic_vector(19 downto 0) := x"0b0a0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_21 : std_logic_vector(19 downto 0) := x"0b0b0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_22 : std_logic_vector(19 downto 0) := x"0b0c0";
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_23 : std_logic_vector(19 downto 0) := x"0b0d0";

  --** FELIG_MON_ITK_STRIPS_ARR
  constant REG_FELIG_MON_ITK_STRIPS_00        : std_logic_vector(19 downto 0) := x"0b0e0";
  constant REG_FELIG_MON_ITK_STRIPS_01        : std_logic_vector(19 downto 0) := x"0b0f0";
  constant REG_FELIG_MON_ITK_STRIPS_02        : std_logic_vector(19 downto 0) := x"0b100";
  constant REG_FELIG_MON_ITK_STRIPS_03        : std_logic_vector(19 downto 0) := x"0b110";
  constant REG_FELIG_MON_ITK_STRIPS_04        : std_logic_vector(19 downto 0) := x"0b120";
  constant REG_FELIG_MON_ITK_STRIPS_05        : std_logic_vector(19 downto 0) := x"0b130";
  constant REG_FELIG_MON_ITK_STRIPS_06        : std_logic_vector(19 downto 0) := x"0b140";
  constant REG_FELIG_MON_ITK_STRIPS_07        : std_logic_vector(19 downto 0) := x"0b150";
  constant REG_FELIG_MON_ITK_STRIPS_08        : std_logic_vector(19 downto 0) := x"0b160";
  constant REG_FELIG_MON_ITK_STRIPS_09        : std_logic_vector(19 downto 0) := x"0b170";
  constant REG_FELIG_MON_ITK_STRIPS_10        : std_logic_vector(19 downto 0) := x"0b180";
  constant REG_FELIG_MON_ITK_STRIPS_11        : std_logic_vector(19 downto 0) := x"0b190";
  constant REG_FELIG_MON_ITK_STRIPS_12        : std_logic_vector(19 downto 0) := x"0b1a0";
  constant REG_FELIG_MON_ITK_STRIPS_13        : std_logic_vector(19 downto 0) := x"0b1b0";
  constant REG_FELIG_MON_ITK_STRIPS_14        : std_logic_vector(19 downto 0) := x"0b1c0";
  constant REG_FELIG_MON_ITK_STRIPS_15        : std_logic_vector(19 downto 0) := x"0b1d0";
  constant REG_FELIG_MON_ITK_STRIPS_16        : std_logic_vector(19 downto 0) := x"0b1e0";
  constant REG_FELIG_MON_ITK_STRIPS_17        : std_logic_vector(19 downto 0) := x"0b1f0";
  constant REG_FELIG_MON_ITK_STRIPS_18        : std_logic_vector(19 downto 0) := x"0b200";
  constant REG_FELIG_MON_ITK_STRIPS_19        : std_logic_vector(19 downto 0) := x"0b210";
  constant REG_FELIG_MON_ITK_STRIPS_20        : std_logic_vector(19 downto 0) := x"0b220";
  constant REG_FELIG_MON_ITK_STRIPS_21        : std_logic_vector(19 downto 0) := x"0b230";
  constant REG_FELIG_MON_ITK_STRIPS_22        : std_logic_vector(19 downto 0) := x"0b240";
  constant REG_FELIG_MON_ITK_STRIPS_23        : std_logic_vector(19 downto 0) := x"0b250";
  constant REG_FMEMU_EVENT_INFO               : std_logic_vector(19 downto 0) := x"0b800";
  constant REG_FMEMU_COUNTERS                 : std_logic_vector(19 downto 0) := x"0b810";
  constant REG_FMEMU_CONTROL                  : std_logic_vector(19 downto 0) := x"0b820";
  constant REG_FMEMU_RANDOM_RAM_ADDR          : std_logic_vector(19 downto 0) := x"0b830";
  constant REG_FMEMU_RANDOM_RAM               : std_logic_vector(19 downto 0) := x"0b840";
  constant REG_FMEMU_RANDOM_CONTROL           : std_logic_vector(19 downto 0) := x"0b850";
  constant REG_FMEMU_CONFIG_WRADDR            : std_logic_vector(19 downto 0) := x"0b860";
  constant REG_FMEMU_CONFIG                   : std_logic_vector(19 downto 0) := x"0b870";

  --** Wishbone
  constant REG_WISHBONE_CONTROL               : std_logic_vector(19 downto 0) := x"0c000";
  constant REG_WISHBONE_WRITE                 : std_logic_vector(19 downto 0) := x"0c010";
  constant REG_WISHBONE_READ                  : std_logic_vector(19 downto 0) := x"0c020";
  constant REG_WISHBONE_STATUS                : std_logic_vector(19 downto 0) := x"0c030";

  --** IPBus
  constant REG_IPBUS_WRITE_ADDRESS            : std_logic_vector(19 downto 0) := x"0c800";
  constant REG_IPBUS_WRITE_DATA               : std_logic_vector(19 downto 0) := x"0c810";
  constant REG_IPBUS_READ_ADDRESS             : std_logic_vector(19 downto 0) := x"0c820";
  constant REG_IPBUS_READ_DATA                : std_logic_vector(19 downto 0) := x"0c830";
  constant REG_IPBUS_PKT_DONE                 : std_logic_vector(19 downto 0) := x"0c840";

  --** ITK_STRIPS_CTRL
  constant REG_GLOBAL_STRIPS_CONFIG           : std_logic_vector(19 downto 0) := x"0d000";
  constant REG_GLOBAL_TRICKLE_TRIGGER         : std_logic_vector(19 downto 0) := x"0d010";
  constant REG_STRIPS_R3_TRIGGER              : std_logic_vector(19 downto 0) := x"0d020";
  constant REG_STRIPS_L1_TRIGGER              : std_logic_vector(19 downto 0) := x"0d030";
  constant REG_STRIPS_R3L1_TRIGGER            : std_logic_vector(19 downto 0) := x"0d040";

  --** MRODregisters
  constant REG_MROD_CTRL                      : std_logic_vector(19 downto 0) := x"0f000";
  constant REG_MROD_TCVRCTRL                  : std_logic_vector(19 downto 0) := x"0f010";
  constant REG_MROD_EP0_CSMENABLE             : std_logic_vector(19 downto 0) := x"0f020";
  constant REG_MROD_EP0_EMPTYSUPPR            : std_logic_vector(19 downto 0) := x"0f030";
  constant REG_MROD_EP0_HPTDCMODE             : std_logic_vector(19 downto 0) := x"0f040";
  constant REG_MROD_EP0_CLRFIFOS              : std_logic_vector(19 downto 0) := x"0f050";
  constant REG_MROD_EP0_EMULOADENA            : std_logic_vector(19 downto 0) := x"0f060";
  constant REG_MROD_EP0_TRXLOOPBACK           : std_logic_vector(19 downto 0) := x"0f070";
  constant REG_MROD_EP0_TXCVRRESET            : std_logic_vector(19 downto 0) := x"0f080";
  constant REG_MROD_EP0_RXRESET               : std_logic_vector(19 downto 0) := x"0f090";
  constant REG_MROD_EP0_TXRESET               : std_logic_vector(19 downto 0) := x"0f0a0";
  constant REG_MROD_EP1_CSMENABLE             : std_logic_vector(19 downto 0) := x"0f0b0";
  constant REG_MROD_EP1_EMPTYSUPPR            : std_logic_vector(19 downto 0) := x"0f0c0";
  constant REG_MROD_EP1_HPTDCMODE             : std_logic_vector(19 downto 0) := x"0f0d0";
  constant REG_MROD_EP1_CLRFIFOS              : std_logic_vector(19 downto 0) := x"0f0e0";
  constant REG_MROD_EP1_EMULOADENA            : std_logic_vector(19 downto 0) := x"0f0f0";
  constant REG_MROD_EP1_TRXLOOPBACK           : std_logic_vector(19 downto 0) := x"0f100";
  constant REG_MROD_EP1_TXCVRRESET            : std_logic_vector(19 downto 0) := x"0f110";
  constant REG_MROD_EP1_RXRESET               : std_logic_vector(19 downto 0) := x"0f120";
  constant REG_MROD_EP1_TXRESET               : std_logic_vector(19 downto 0) := x"0f130";

  --** MRODmonitors
  constant REG_MROD_EP0_CSMH_EMPTY            : std_logic_vector(19 downto 0) := x"0f800";
  constant REG_MROD_EP0_CSMH_FULL             : std_logic_vector(19 downto 0) := x"0f810";
  constant REG_MROD_EP0_RXALIGNBSY            : std_logic_vector(19 downto 0) := x"0f820";
  constant REG_MROD_EP0_RXRECDATA             : std_logic_vector(19 downto 0) := x"0f830";
  constant REG_MROD_EP0_RXRECIDLES            : std_logic_vector(19 downto 0) := x"0f840";
  constant REG_MROD_EP0_TXLOCKED              : std_logic_vector(19 downto 0) := x"0f850";
  constant REG_MROD_EP1_CSMH_EMPTY            : std_logic_vector(19 downto 0) := x"0f860";
  constant REG_MROD_EP1_CSMH_FULL             : std_logic_vector(19 downto 0) := x"0f870";
  constant REG_MROD_EP1_RXALIGNBSY            : std_logic_vector(19 downto 0) := x"0f880";
  constant REG_MROD_EP1_RXRECDATA             : std_logic_vector(19 downto 0) := x"0f890";
  constant REG_MROD_EP1_RXRECIDLES            : std_logic_vector(19 downto 0) := x"0f8a0";
  constant REG_MROD_EP1_TXLOCKED              : std_logic_vector(19 downto 0) := x"0f8b0";
  -----------------------------------
  ---- GENERATED code END #1 ##  ----
  -----------------------------------

  --!
  --! --> CONTROL: Read/Write User Application Registers (Written by PCIe)
  ------------------------------------
  ---- ## GENERATED code BEGIN #2 ----
  ------------------------------------
  -- Bitfields of Control Record
  type bitfield_timeout_ctrl_w_type is record
    ENABLE                         : std_logic_vector(32 downto 32);  -- 1 enables the timout trailer generation for ToHost mode
    TIMEOUT                        : std_logic_vector(31 downto 0);   -- Number of 40 MHz clock cycles after which a timeout occurs.
  end record;

  type bitfield_crtohost_fifo_status_t_type is record
    CLEAR                          : std_logic_vector(64 downto 64);  -- Any write to this register clears the latched FULL flags
  end record;

  type bitfield_crtohost_dma_descriptor_1_t_type is record
    WR_EN                          : std_logic_vector(64 downto 64);  -- Any write to this register assigns the DMA ID to the AXIS_ID set in CRTOHOST_DMA_DESCRIPTOR_2.AXIS_ID
    DESCR                          : std_logic_vector(2 downto 0);    -- Target descriptor
  end record;

  type bitfield_crtohost_dma_descriptor_2_w_type is record
    AXIS_ID                        : std_logic_vector(10 downto 0);   -- ID of the AXI stream (E-Path ID) to associate with CRTOHOST_DMA_DESCRIPTOR_1.DESCR
  end record;

  type bitfield_crfromhost_fifo_status_t_type is record
    CLEAR                          : std_logic_vector(64 downto 64);  -- Any write to this register clears the latched FULL flags
  end record;

  --Array of registers (std_logic_vector)
  type bitfield_broadcast_enable_w_array_type is  array (0 to 23) of  std_logic_vector(41 downto 0);   -- Enable path to be included in a broadcast message.
  type bitfield_has_stream_id_w_type is record
    EGROUP6                        : std_logic_vector(55 downto 48);  -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
    EGROUP5                        : std_logic_vector(47 downto 40);  -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
    EGROUP4                        : std_logic_vector(39 downto 32);  -- EPATH is associated with a STREAM ID
    EGROUP3                        : std_logic_vector(31 downto 24);  -- EPATH is associated with a STREAM ID
    EGROUP2                        : std_logic_vector(23 downto 16);  -- EPATH is associated with a STREAM ID
    EGROUP1                        : std_logic_vector(15 downto 8);   -- EPATH is associated with a STREAM ID
    EGROUP0                        : std_logic_vector(7 downto 0);    -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  end record;
  --Array of registers
  type bitfield_has_stream_id_w_array_type is array (0 to 23) of bitfield_has_stream_id_w_type;
  type bitfield_decoding_egroup_ctrl_w_type is record
    ENABLE_TRUNCATION              : std_logic_vector(59 downto 59);  -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
    REVERSE_ELINKS                 : std_logic_vector(50 downto 43);  -- enables bit reversing for the elink in the given epath
    PATH_ENCODING                  : std_logic_vector(42 downto 11);  -- Encoding for every EPATH, 4 bits per E-path
                                                                      -- 0: direct mode
                                                                      -- 1: 8b10b mode
                                                                      -- 2: HDLC mode
                                                                      -- 3: TTC
                                                                      -- 4: ITk Strips 8b10b
                                                                      -- 5: ITk Pixel
                                                                      -- 6: Endeavour
                                                                      -- 7-15:  reserved
                                                                      
    EPATH_WIDTH                    : std_logic_vector(10 downto 8);   -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
    EPATH_ENA                      : std_logic_vector(7 downto 0);    -- Enable bits per EPATH
  end record;
  --Array of registers
  type bitfield_decoding_egroup_ctrl_w_array_type is array (0 to 6) of bitfield_decoding_egroup_ctrl_w_type;
  --Two dimensional array of registers
  type bitfield_decoding_egroup_ctrl_w_2d_array_type is array (0 to 11) of bitfield_decoding_egroup_ctrl_w_array_type;
  type bitfield_mini_egroup_tohost_w_type is record
    ENABLE_AUX_TRUNCATION          : std_logic_vector(15 downto 15);  -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
    ENABLE_IC_TRUNCATION           : std_logic_vector(14 downto 14);  -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
    ENABLE_EC_TRUNCATION           : std_logic_vector(13 downto 13);  -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
    AUX_BIT_SWAPPING               : std_logic_vector(11 downto 11);  -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
    AUX_ENABLE                     : std_logic_vector(10 downto 10);  -- Enables the AUX channel
    IC_BIT_SWAPPING                : std_logic_vector(8 downto 8);    -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
    IC_ENABLE                      : std_logic_vector(7 downto 7);    -- Enables the IC channel
    EC_BIT_SWAPPING                : std_logic_vector(5 downto 5);    -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
    EC_ENCODING                    : std_logic_vector(4 downto 1);    -- Configures encoding of the EC channel
    EC_ENABLE                      : std_logic_vector(0 downto 0);    -- Enables the EC channel
  end record;
  --Array of registers
  type bitfield_mini_egroup_tohost_w_array_type is array (0 to 23) of bitfield_mini_egroup_tohost_w_type;
  type bitfield_yarr_debug_allegroup_tohost_w_type is record
    REF_PACKET                     : std_logic_vector(63 downto 32);  -- Reference packet to be matched
  end record;
  --Array of registers
  type bitfield_yarr_debug_allegroup_tohost_w_array_type is array (0 to 11) of bitfield_yarr_debug_allegroup_tohost_w_type;
  --Array of registers (std_logic_vector)
  type bitfield_super_chunk_factor_link_w_array_type is  array (0 to 11) of  std_logic_vector(7 downto 0);    -- number of chunks glued together
  type bitfield_decoding_link_cb_w_type is record
    CBOPT                          : std_logic_vector(3 downto 0);    -- Channel bonding option
                                                                      -- 0: no bonding
                                                                      -- 3: Bonding 0/1/2 3/4/5
                                                                      -- other values: reserved
                                                                      
  end record;
  --Array of registers
  type bitfield_decoding_link_cb_w_array_type is array (0 to 11) of bitfield_decoding_link_cb_w_type;
  type bitfield_encoding_egroup_ctrl_w_type is record
    ENABLE_DELAY                   : std_logic_vector(63 downto 63);  -- Enable inter-packet delay generation in HDLC encoder
    TTC_OPTION                     : std_logic_vector(62 downto 59);  -- Selects TTC bits sent to the E-link
    REVERSE_ELINKS                 : std_logic_vector(50 downto 43);  -- enables bit reversing for the elink in the given epath
    EPATH_WIDTH                    : std_logic_vector(42 downto 40);  -- Width of the Elinks in the egroup
                                                                      -- 0: 2 bit 80 Mb/s
                                                                      -- 1: 4 bit 160 Mb/s
                                                                      -- 2: 8 bit 320 Mb/s
                                                                      
    PATH_ENCODING                  : std_logic_vector(39 downto 8);   -- Encoding for every EPATH, 4 bits per E-Path
                                                                      -- 0: No encoding
                                                                      -- 1: 8b10b mode
                                                                      -- 2: HDLC mode
                                                                      -- 3: ITk Strip LCB
                                                                      -- 4: ITk Pixel
                                                                      -- 5: Endeavour
                                                                      -- 6: reserved
                                                                      -- 7: reserved
                                                                      -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                      
    EPATH_ENA                      : std_logic_vector(7 downto 0);    -- Enable bits per E-PATH
  end record;
  --Array of registers
  type bitfield_encoding_egroup_ctrl_w_array_type is array (0 to 4) of bitfield_encoding_egroup_ctrl_w_type;
  --Two dimensional array of registers
  type bitfield_encoding_egroup_ctrl_w_2d_array_type is array (0 to 11) of bitfield_encoding_egroup_ctrl_w_array_type;
  type bitfield_mini_egroup_fromhost_w_type is record
    ENABLE_DELAY                   : std_logic_vector(13 downto 13);  -- Enable inter-packet delay generation in HDLC encoder
    AUX_BIT_SWAPPING               : std_logic_vector(11 downto 11);  -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
    AUX_ENABLE                     : std_logic_vector(10 downto 10);  -- Enables the AUX channel
    IC_BIT_SWAPPING                : std_logic_vector(8 downto 8);    -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
    IC_ENABLE                      : std_logic_vector(7 downto 7);    -- Enables the IC channel
    EC_BIT_SWAPPING                : std_logic_vector(5 downto 5);    -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
    EC_ENCODING                    : std_logic_vector(4 downto 1);    -- Configures encoding of the EC channel
    EC_ENABLE                      : std_logic_vector(0 downto 0);    -- Configures the FromHost Mini egroup
  end record;
  --Array of registers
  type bitfield_mini_egroup_fromhost_w_array_type is array (0 to 23) of bitfield_mini_egroup_fromhost_w_type;
  type bitfield_encoding_egroup_fei4_ctrl_w_type is record
    PHASE_DELAY1                   : std_logic_vector(11 downto 9);   -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
    MANCHESTER_ENABLE1             : std_logic_vector(8 downto 8);    -- enable manchester encoding
    AUTOMATIC_MERGE_DISABLE1       : std_logic_vector(7 downto 7);    -- Disable automatic merging
    TTC_SELECT1                    : std_logic_vector(6 downto 6);    -- TTC/FromHost select (if automatic merging is disabled)
    PHASE_DELAY0                   : std_logic_vector(5 downto 3);    -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
    MANCHESTER_ENABLE0             : std_logic_vector(2 downto 2);    -- enable manchester encoding
    AUTOMATIC_MERGE_DISABLE0       : std_logic_vector(1 downto 1);    -- Disable automatic merging
    TTC_SELECT0                    : std_logic_vector(0 downto 0);    -- TTC/FromHost select (if automatic merging is disabled)
  end record;
  --Array of registers
  type bitfield_encoding_egroup_fei4_ctrl_w_array_type is array (0 to 4) of bitfield_encoding_egroup_fei4_ctrl_w_type;
  --Two dimensional array of registers
  type bitfield_encoding_egroup_fei4_ctrl_w_2d_array_type is array (0 to 11) of bitfield_encoding_egroup_fei4_ctrl_w_array_type;
  type bitfield_yarr_debug_allegroup_fromhost1_w_type is record
    RD53A_AZ_EN                    : std_logic_vector(48 downto 48);  -- Auto zeroing module enable
    REF_DLY_GENCALTRIG             : std_logic_vector(7 downto 0);    -- Reference distance between GenCal and First Trigger
  end record;
  --Array of registers
  type bitfield_yarr_debug_allegroup_fromhost1_w_array_type is array (0 to 11) of bitfield_yarr_debug_allegroup_fromhost1_w_type;
  type bitfield_yarr_debug_allegroup_fromhost2_w_type is record
    REF_CMD                        : std_logic_vector(15 downto 0);   -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  end record;
  --Array of registers
  type bitfield_yarr_debug_allegroup_fromhost2_w_array_type is array (0 to 11) of bitfield_yarr_debug_allegroup_fromhost2_w_type;
  type bitfield_fe_emu_ena_w_type is record
    EMU_TOFRONTEND                 : std_logic_vector(1 downto 1);    -- Enable GBT dummy emulator ToFrontEnd
    EMU_TOHOST                     : std_logic_vector(0 downto 0);    -- Enable GBT dummy emulator ToHost
  end record;

  type bitfield_fe_emu_config_w_type is record
    WE                             : std_logic_vector(54 downto 47);  -- write enable array, every bit is one emulator RAM block
    WRADDR                         : std_logic_vector(46 downto 33);  -- write address bus
    WRDATA                         : std_logic_vector(32 downto 0);   -- write data bus
  end record;

  type bitfield_fe_emu_read_w_type is record
    SEL                            : std_logic_vector(35 downto 33);  -- Select ramblock to read back
  end record;

  type bitfield_fe_emu_logic_w_type is record
    L1A_TRIGGERED                  : std_logic_vector(33 downto 33);  -- 1 Send a chunk on every L1A, 0 use the IDLES to determine the rate
    ENA                            : std_logic_vector(32 downto 32);  -- Enable logic based FrontEnd emulator, instead of RAM based.
    IDLES                          : std_logic_vector(31 downto 16);  -- Number of IDLE bytes between chunks.
    CHUNK_LENGTH                   : std_logic_vector(15 downto 0);   -- Chunk length in bytes
  end record;

  type bitfield_gbt_mode_ctrl_w_type is record
    RX_ALIGN_TB_SW                 : std_logic_vector(2 downto 2);    -- RX_ALIGN_TB_SW
    RX_ALIGN_SW                    : std_logic_vector(1 downto 1);    -- RX_ALIGN_SW
    DESMUX_USE_SW                  : std_logic_vector(0 downto 0);    -- DESMUX_USE_SW
  end record;

  type bitfield_gbt_pll_reset_w_type is record
    QPLL_RESET                     : std_logic_vector(59 downto 48);  -- QPLL_RESET [11:0]
    CPLL_RESET                     : std_logic_vector(47 downto 0);   -- CPLL_RESET [47:0]
  end record;

  type bitfield_gbt_soft_tx_reset_w_type is record
    RESET_ALL                      : std_logic_vector(59 downto 48);  -- SOFT_TX_RESET_ALL [11:0]
    RESET_GT                       : std_logic_vector(47 downto 0);   -- SOFT_TX_RESET_GT [47:0]
  end record;

  type bitfield_gbt_soft_rx_reset_w_type is record
    RESET_ALL                      : std_logic_vector(59 downto 48);  -- SOFT_TX_RESET_ALL [11:0]
    RESET_GT                       : std_logic_vector(47 downto 0);   -- SOFT_TX_RESET_GT [47:0]
  end record;

  type bitfield_gbt_tohost_fanout_w_type is record
    LOCK                           : std_logic_vector(48 downto 48);  -- Locks this particular register. If set prevents software from touching it.
    SEL                            : std_logic_vector(47 downto 0);   -- ToHost FanOut/Selector. Every bitfield is a channel:
                                                                      --   1 : GBT_EMU, select GBT Emulator for a specific CentralRouter channel
                                                                      --   0 : GBT_WRAP, select real GBT link for a specific CentralRouter channel
                                                                      
  end record;

  type bitfield_gbt_tofrontend_fanout_w_type is record
    LOCK                           : std_logic_vector(48 downto 48);  -- Locks this particular register. If set prevents software from touching it.
    SEL                            : std_logic_vector(47 downto 0);   -- ToFrontEnd FanOut/Selector. Every bitfield is a channel:
                                                                      --   1 : GBT_EMU, select GBT Emulator for a specific GBT link
                                                                      --   0 : TTC_DEC, select CentralRouter data (including TTC) for a specific GBT link
                                                                      --   
                                                                      
  end record;

  type bitfield_fullmode_auto_rx_reset_w_type is record
    ENABLE                         : std_logic_vector(32 downto 32);  -- Enable the Automatic RX Reset mechanism
    TIMEOUT                        : std_logic_vector(31 downto 0);   -- Number of 40 MHz clock cycles until an unaligned link results in a reset pulse
  end record;

  type bitfield_ttc_dec_ctrl_w_type is record
    B_CHAN_DELAY                   : std_logic_vector(30 downto 27);  -- Number of BC to delay the L1A distribution to the frontends
    BCID_ONBCR                     : std_logic_vector(26 downto 15);  -- BCID is set to this value when BCR arrives
    ECR_BCR_SWAP                   : std_logic_vector(13 downto 13);  -- ECR and BCR signals are swapped at the output of the TTC decoder (needed only for LAr TTC)
    BUSY_OUTPUT_INHIBIT            : std_logic_vector(12 downto 12);  -- forces the Busy LEMO output to BUSY-OFF
    TOHOST_RST                     : std_logic_vector(11 downto 11);  -- reset toHost in ttc decoder
    TT_BCH_EN                      : std_logic_vector(10 downto 10);  -- trigger type enable / disable for TTC-ToHost
    XL1ID_SW                       : std_logic_vector(9 downto 2);    -- set XL1ID value, the value to be set by XL1ID_RST signal
    XL1ID_RST                      : std_logic_vector(1 downto 1);    -- giving a trigger signal to reset XL1ID value
    MASTER_BUSY                    : std_logic_vector(0 downto 0);    -- L1A trigger throttling
  end record;

  type bitfield_ttc_emu_w_type is record
    SEL                            : std_logic_vector(1 downto 1);    -- Select TTC data source 1 TTC Emu | 0 TTC Decoder
    ENA                            : std_logic_vector(0 downto 0);    -- Clear to load into the TTC emulator’s memory the required sequence, Set to run the TTC emulator sequence
  end record;

  type bitfield_ttc_busy_timing_ctrl_w_type is record
    PRESCALE                       : std_logic_vector(51 downto 32);  -- Prescales the 40MHz clock to create an internal slow clock
    BUSY_WIDTH                     : std_logic_vector(31 downto 16);  -- Minimum number of 40MHz clocks that the busy is asserted
    LIMIT_TIME                     : std_logic_vector(15 downto 0);   -- Number of prescaled clocks a given busy must be asserted before it is recognized
  end record;

  type bitfield_ttc_emu_control_w_type is record
    BUSY_IN_ENABLE                 : std_logic_vector(33 downto 33);  -- Enable internal BUSY input to stop L1A on BUSY
    BROADCAST                      : std_logic_vector(32 downto 27);  -- Broadcast data
    ECR                            : std_logic_vector(26 downto 26);  -- Event counter reset
    BCR                            : std_logic_vector(25 downto 25);  -- Bunch counter reset
    L1A                            : std_logic_vector(24 downto 24);  -- Level 1 Accept
  end record;

  type bitfield_ttc_ecr_monitor_t_type is record
    CLEAR                          : std_logic_vector(64 downto 64);  -- Counts the number of ECRs received from the TTC system, any write to this register clears the counter
  end record;

  type bitfield_ttc_ttype_monitor_t_type is record
    CLEAR                          : std_logic_vector(64 downto 64);  -- Counts the number of TType received from the TTC system, any write to this register clears the counter
  end record;

  type bitfield_ttc_bcr_periodicity_monitor_t_type is record
    CLEAR                          : std_logic_vector(64 downto 64);  -- Counts the number of times the BCR period does not match 3564, any write to this register clears the counter
  end record;

  type bitfield_ttc_bcr_counter_t_type is record
    CLEAR                          : std_logic_vector(64 downto 64);  -- Counts the number of times BCR is issued, any write to this register clears the counter
  end record;

  type bitfield_xoff_fm_high_thresh_t_type is record
    CLEAR_LATCH                    : std_logic_vector(64 downto 64);  -- Writing this register will clear all CROSS_LATCHED bits
  end record;

  type bitfield_dma_busy_status_t_type is record
    CLEAR_LATCH                    : std_logic_vector(64 downto 64);  -- Any write to this register clears TOHOST_BUSY_LATCHED
    ENABLE                         : std_logic_vector(4 downto 4);    -- Enable the DMA buffer on the server as a source of busy
  end record;

  type bitfield_fm_busy_channel_status_t_type is record
    CLEAR_LATCH                    : std_logic_vector(64 downto 64);  -- Any write to this register will clear the BUSY_LATCHED bits
  end record;

  type bitfield_busy_main_output_fifo_thresh_w_type is record
    BUSY_ENABLE                    : std_logic_vector(24 downto 24);  -- Enable busy generation if thresholds are crossed
    LOW                            : std_logic_vector(23 downto 12);  -- Low, Negate threshold of busy generation from main output fifo
    HIGH                           : std_logic_vector(11 downto 0);   -- High, Assert threshold of busy generation from main output fifo
  end record;

  type bitfield_busy_main_output_fifo_status_t_type is record
    CLEAR_LATCHED                  : std_logic_vector(64 downto 64);  -- Any write to this register will clear the
  end record;

  --Array of registers (std_logic_vector)
  type bitfield_elink_busy_enable_w_array_type is  array (0 to 23) of  std_logic_vector(56 downto 0);   -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  type bitfield_hk_ctrl_i2c_w_type is record
    CONFIG_TRIG                    : std_logic_vector(1 downto 1);    -- i2c_config_trig
    CLKFREQ_SEL                    : std_logic_vector(0 downto 0);    -- i2c_clkfreq_sel
  end record;

  type bitfield_hk_ctrl_fmc_w_type is record
    SI5345_INSEL                   : std_logic_vector(6 downto 5);    -- Selects the input clock source
                                                                      --   0 : FPGA (FMC LA01)
                                                                      --   1 : FMC OSC (40.079 MHz)
                                                                      --   2 : FPGA (FMC LA18)
                                                                      
    SI5345_A                       : std_logic_vector(4 downto 3);    -- Si5345 I2C address select 2 LSB (0x0:default, dev id 0x68)
    SI5345_OE                      : std_logic_vector(2 downto 2);    -- Si5345 active low output enable  (0:enable)
    SI5345_RSTN                    : std_logic_vector(1 downto 1);    -- Si5345 active low output enable  (0:reset)
    SI5345_SEL                     : std_logic_vector(0 downto 0);    -- Si5345 programming mode
                                                                      --   1 : I2C mode (default)
                                                                      --   0 : SPI mode
                                                                      
  end record;

  type bitfield_hk_mon_fmc_w_type is record
    SI5345_LOL                     : std_logic_vector(1 downto 1);    -- Si5345 Loss Of Lock pin
    SI5345_INTR                    : std_logic_vector(0 downto 0);    -- Si5345 Interrupt flagging chip change of status
  end record;

  type bitfield_mmcm_main_w_type is record
    LCLK_SEL                       : std_logic_vector(3 downto 3);    -- 1: LCLK
                                                                      -- 0: TTC
                                                                      
  end record;

  type bitfield_i2c_wr_t_type is record
    I2C_WREN                       : std_logic_vector(64 downto 64);  -- Any write to this register triggers an I2C read or write sequence
    WRITE_2BYTES                   : std_logic_vector(24 downto 24);  -- Write two bytes
    DATA_BYTE2                     : std_logic_vector(23 downto 16);  -- Data byte 2
    DATA_BYTE1                     : std_logic_vector(15 downto 8);   -- Data byte 1
    SLAVE_ADDRESS                  : std_logic_vector(7 downto 1);    -- Slave address
    READ_NOT_WRITE                 : std_logic_vector(0 downto 0);    -- READ/<o>WRITE</o>
  end record;

  type bitfield_i2c_rd_t_type is record
    I2C_RDEN                       : std_logic_vector(64 downto 64);  -- Any write to this register pops the last I2C data from the FIFO
  end record;

  type bitfield_int_test_t_type is record
    TRIGGER                        : std_logic_vector(64 downto 64);  -- Fire a test MSIx interrupt set in IRQ
    IRQ                            : std_logic_vector(3 downto 0);    -- Set this field to a value equal to the MSIX interrupt to be fired. The write triggers the interrupt immediately.
  end record;

  type bitfield_config_flash_wr_w_type is record
    FAST_WRITE                     : std_logic_vector(57 downto 57);  -- Write command only. Only used for fast programming.
    FAST_READ                      : std_logic_vector(56 downto 56);  -- Status reading without command writing. Only used for fast programming.
    PAR_CTRL                       : std_logic_vector(55 downto 55);  -- Choose use FW or uC to select the Flash partition. 1 FW | 0 uC.
    PAR_WR                         : std_logic_vector(54 downto 53);  -- Choose Flash partition. Valid when PAR_CTRL is 1.
    FLASH_SEL                      : std_logic_vector(52 downto 52);  -- 1 takes control over flash, 0 gives JTAG control over flash
    DO_INIT                        : std_logic_vector(51 downto 51);  -- Untested feature, don't use it yet.
    DO_READSTATUS                  : std_logic_vector(50 downto 50);  -- Reads status from flash
    DO_CLEARSTATUS                 : std_logic_vector(49 downto 49);  -- Clears status reading from flash, back to normal flash operation
    DO_ERASEBLOCK                  : std_logic_vector(48 downto 48);  -- Erased the current block of the flash, this register has to be cleared by software
    DO_UNLOCK_BLOCK                : std_logic_vector(47 downto 47);  -- Unlock writes to the current block, this register has to be cleared by software
    DO_READ                        : std_logic_vector(46 downto 46);  -- Reads the 16 bits from current address, this register has to be cleared by software
    DO_WRITE                       : std_logic_vector(45 downto 45);  -- Writes the 16 bits to current address, this register has to be cleared by software
    DO_READDEVICEID                : std_logic_vector(44 downto 44);  -- DIN should return 0x0089, this register has to be cleared by software
    DO_RESET                       : std_logic_vector(43 downto 43);  -- Can be used in the future, currently disconnected in firmware
    ADDRESS                        : std_logic_vector(42 downto 16);  -- Address for read and write operations (25 bits, upper 2 bits are controlled by uC)
    WRITE_DATA                     : std_logic_vector(15 downto 0);   -- Value of data to write towards flash
  end record;

  type bitfield_rxusrclk_freq_w_type is record
    CHANNEL                        : std_logic_vector(37 downto 32);  -- Select the Transceiver channel to measure the clock from.
  end record;

  type bitfield_felig_data_gen_config_w_type is record
    USERDATA                       : std_logic_vector(63 downto 48);  -- Sets static payload word. When PATTERN_SEL=1.
    CHUNK_LENGTH                   : std_logic_vector(47 downto 32);  -- FELIG data generator chunk-length in bytes.
    RESET                          : std_logic_vector(19 downto 15);  -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
    SW_BUSY                        : std_logic_vector(14 downto 10);  -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
    DATA_FORMAT                    : std_logic_vector(9 downto 5);    -- FELIG data generator format. 0:8b10b, 1:direct.
    PATTERN_SEL                    : std_logic_vector(4 downto 0);    -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  end record;
  --Array of registers
  type bitfield_felig_data_gen_config_w_array_type is array (0 to 23) of bitfield_felig_data_gen_config_w_type;
  type bitfield_felig_elink_config_w_type is record
    ENDIAN_MOD                     : std_logic_vector(39 downto 35);  -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
    INPUT_WIDTH                    : std_logic_vector(34 downto 30);  -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
    OUTPUT_WIDTH                   : std_logic_vector(9 downto 0);    -- FELIG elink data output width.
  end record;
  --Array of registers
  type bitfield_felig_elink_config_w_array_type is array (0 to 23) of bitfield_felig_elink_config_w_type;
  --Array of registers (std_logic_vector)
  type bitfield_felig_elink_enable_w_array_type is  array (0 to 23) of  std_logic_vector(39 downto 0);   -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  type bitfield_felig_global_control_w_type is record
    FAKE_L1A_RATE                  : std_logic_vector(63 downto 36);  -- Sets the internal fake L1 trigger rate. [25ns/LSB]
    PICXO_OFFSET_PPM               : std_logic_vector(35 downto 14);  -- When OFFSET_EN is 1, this directly sets the output frequency, within the given adjustment range.
    TRACK_DATA                     : std_logic_vector(12 downto 12);  -- FELIG GT core control.  Must be set to enable normal operation.
    RXUSERRDY                      : std_logic_vector(11 downto 11);  -- FELIG GT core control.  Must be set to enable normal operation.
    TXUSERRDY                      : std_logic_vector(10 downto 10);  -- FELIG GT core control.  Must be set to enable normal operation.
    AUTO_RESET                     : std_logic_vector(9 downto 9);    -- FELIG GT core control.  If set the GT core automatically resets on data error.
    PICXO_RESET                    : std_logic_vector(8 downto 8);    -- FELIG GT core control.  Manual PICXO reset.
    GTTX_RESET                     : std_logic_vector(7 downto 7);    -- FELIG GT core control.  Manual GT TX reset
    CPLL_RESET                     : std_logic_vector(6 downto 6);    -- FELIG GT core control.  Manual CPLL reset.
    X3_X4_OUTPUT_SELECT            : std_logic_vector(5 downto 0);    -- X3/X4 SMA output source select.
  end record;

  type bitfield_felig_lane_config_w_type is record
    B_CH_BIT_SEL                   : std_logic_vector(63 downto 42);  -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
    A_CH_BIT_SEL                   : std_logic_vector(41 downto 35);  -- Selects the bit from the received FELIX data from which to extract the L1A.
    LB_FIFO_DELAY                  : std_logic_vector(34 downto 30);  -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
    ELINK_SYNC                     : std_logic_vector(7 downto 7);    -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
    PICXO_OFFEST_EN                : std_logic_vector(6 downto 6);    -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
    PI_HOLD                        : std_logic_vector(5 downto 5);    -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
    GBT_LB_ENABLE                  : std_logic_vector(4 downto 4);    -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
    GBH_LB_ENABLE                  : std_logic_vector(3 downto 3);    -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
    L1A_SOURCE                     : std_logic_vector(2 downto 2);    -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
    GBT_EMU_SOURCE                 : std_logic_vector(1 downto 1);    -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
    FG_SOURCE                      : std_logic_vector(0 downto 0);    -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  end record;
  --Array of registers
  type bitfield_felig_lane_config_w_array_type is array (0 to 23) of bitfield_felig_lane_config_w_type;
  type bitfield_felig_mon_freq_global_w_type is record
    XTAL_100MHZ                    : std_logic_vector(63 downto 32);  -- FELIG local oscillator frequency[Hz].
    CLK_41_667MHZ                  : std_logic_vector(31 downto 0);   -- FELIG PCIE MGTREFCLK frequency[Hz].
  end record;

  type bitfield_felig_reset_w_type is record
    LB_FIFO                        : std_logic_vector(63 downto 48);  -- One bit per lane.  When set to 1, resets all loopback FIFOs.
    FRAMEGEN                       : std_logic_vector(47 downto 24);  -- One bit per lane.  When set to 1, resets all FELIG link checking logic.
    LANE                           : std_logic_vector(23 downto 0);   -- One bit per lane.  When set to 1, resets all FELIG lane logic.
  end record;

  type bitfield_felig_itk_strips_data_gen_config_w_type is record
    ITKS_FIFO_CTL                  : std_logic_vector(19 downto 17);  -- data fifo control 2:rst 1:rd 0:wr.
    ITKS_FIFO_DATA                 : std_logic_vector(16 downto 0);   -- itks emu data 16:last word 15-0:data word
  end record;
  --Array of registers
  type bitfield_felig_itk_strips_data_gen_config_w_array_type is array (0 to 23) of bitfield_felig_itk_strips_data_gen_config_w_type;
  type bitfield_fmemu_counters_w_type is record
    WORD_CNT                       : std_logic_vector(63 downto 48);  -- Number of 32b words in one chunk
    IDLE_CNT                       : std_logic_vector(47 downto 32);  -- Minimum number of idles between chunks
    L1A_CNT                        : std_logic_vector(31 downto 16);  -- Number of chunks to send if not in TTC mode
    BUSY_TH_HIGH                   : std_logic_vector(15 downto 8);   -- Assert BUSY-ON above this threshold
    BUSY_TH_LOW                    : std_logic_vector(7 downto 0);    -- De-assert BUSY-ON below this threshold
  end record;

  type bitfield_fmemu_control_w_type is record
    L1A_BITNR                      : std_logic_vector(63 downto 56);  -- Bitfield for L1A in TTC frame
    XONXOFF_BITNR                  : std_logic_vector(55 downto 48);  -- Bitfield for Xon/Xoff in TTC frame
    EMU_START                      : std_logic_vector(47 downto 47);  -- Start emulator functionality
    TTC_MODE                       : std_logic_vector(46 downto 46);  -- Control the emulator by TTC input or by RegMap (1/0)
    XONXOFF                        : std_logic_vector(45 downto 45);  -- Enable Xon/Xoff functionality (1/0)
    INLC_CRC32                     : std_logic_vector(44 downto 44);  -- 0: No checksum
                                                                      -- 1: Append the data with a CRC32
                                                                      
    BCR                            : std_logic_vector(43 downto 43);  -- Reset BCID to 0
    ECR                            : std_logic_vector(42 downto 42);  -- Reset L1ID to 0
    CONSTANT_CHUNK_LENGTH          : std_logic_vector(41 downto 41);  -- Data source select
                                                                      -- 0: Random chunk length
                                                                      -- 1: Constant chunk length
                                                                      
    FFU_FM_EMU_T                   : std_logic_vector(16 downto 16);  -- For Future Use (trigger registers)
    FE_BUSY_ENABLE                 : std_logic_vector(0 downto 0);    -- Enable the BUSY mechanism if L1A counter passes threshold
  end record;

  type bitfield_fmemu_random_ram_t_type is record
    WE                             : std_logic_vector(64 downto 64);  -- Any write to this register (DATA) triggers a write to the ramblock
    CHANNEL_SELECT                 : std_logic_vector(39 downto 16);  -- Enable write enable only for the selected channel
    DATA                           : std_logic_vector(15 downto 0);   -- DATA field to be written to FMEMU_RANDOM_RAM_ADDR
  end record;

  type bitfield_fmemu_random_control_w_type is record
    SELECT_RANDOM                  : std_logic_vector(20 downto 20);  -- 1 enables the random chunk length, 0 uses a constant chunk length
    SEED                           : std_logic_vector(19 downto 10);  -- Seed for the random number generator, should not be 0
    POLYNOMIAL                     : std_logic_vector(9 downto 0);    -- POLYNOMIAL for the random number generator (10b LFSR) Bit9 should always be 1
  end record;

  type bitfield_fmemu_config_t_type is record
    WE                             : std_logic_vector(64 downto 64);  -- Any write to register WRDATA triggers a write to the ramblock
    CHANNEL_SELECT                 : std_logic_vector(55 downto 32);  -- Enable write enable only for the selected channel
    WRDATA                         : std_logic_vector(31 downto 0);   -- DATA field to be written to FMEMU_RANDOM_RAM_ADDR
  end record;

  type bitfield_wishbone_control_w_type is record
    WRITE_NOT_READ                 : std_logic_vector(32 downto 32);  -- wishbone write command wishbone read command
    ADDRESS                        : std_logic_vector(31 downto 0);   -- Slave address for Wishbone bus
  end record;

  type bitfield_wishbone_write_t_type is record
    WRITE_ENABLE                   : std_logic_vector(64 downto 64);  -- Any write to this register triggers a write to the Wupper to Wishbone fifo
    DATA                           : std_logic_vector(31 downto 0);   -- Wishbone
  end record;

  type bitfield_wishbone_read_t_type is record
    READ_ENABLE                    : std_logic_vector(64 downto 64);  -- Any write to this register triggers a read from the Wishbone to Wupper fifo
  end record;

  type bitfield_ipbus_write_data_t_type is record
    WRITE_ENABLE                   : std_logic_vector(64 downto 64);  -- Any write to this register triggers a write to the Wupper to IPBus inout RAM
    DATA                           : std_logic_vector(63 downto 0);   -- IPbus data to write to RAM
  end record;

  type bitfield_global_strips_config_w_type is record
    TEST_MODULE_MASK               : std_logic_vector(63 downto 59);  -- (for tests only) contains R3 mask for the simulated trigger data
    TEST_R3L1_TAG                  : std_logic_vector(58 downto 52);  -- (for tests only) contains R3 or L1 tag for the simulated trigger data
    TTC_GENERATE_GATING_ENABLE     : std_logic_vector(51 downto 51);  -- Global control for gating signal generation. Enables generating trickle gating signal in response to TTC BCR. TRICKLE_TRIG_RUN must also be enabled for the trickle configuration to work. (See also BC_START, and BC_STOP fields)
    TTC_GATING_OVERRIDE            : std_logic_vector(50 downto 50);  -- Overrides and disables gating signal generation when set to '1' (use if the elink is deadlocked and commands don't reach it).
    INVERT_AMAC_IN                 : std_logic_vector(4 downto 4);    -- Invert the polarity of all FELIX AMAC_IN elinks
    INVERT_AMAC_OUT                : std_logic_vector(3 downto 3);    -- Invert the polarity of all FELIX AMAC_OUT elinks
    INVERT_DIN                     : std_logic_vector(2 downto 2);    -- Invert the polarity of all FELIX 8-bit IN 8b10b elinks
    INVERT_R3L1_OUT                : std_logic_vector(1 downto 1);    -- Invert the polarity of all FELIX R3L1 elinks
    INVERT_LCB_OUT                 : std_logic_vector(0 downto 0);    -- Invert the polarity of all FELIX LCB elinks
  end record;

  type bitfield_mrod_ctrl_w_type is record
    OPTIONS                        : std_logic_vector(15 downto 8);   -- Extra options for MROD
    ENASPARE1                      : std_logic_vector(7 downto 7);    -- Enable spare1
    ENAMANSLIDE                    : std_logic_vector(6 downto 6);    -- Enable Manual Slide in Rx Locking
    ENAPASSALL                     : std_logic_vector(5 downto 5);    -- Enable PassAll in EmptySuppress
    ENATXCOUNT                     : std_logic_vector(4 downto 4);    -- Enable SimpleCount in TxDriver for locking
    GOLTESTMODE                    : std_logic_vector(3 downto 0);    -- GOL Test Mode (emulate CSM):
                                                                      --   0: Run Data Emulator when 1;     0: stop, load emulator fifo
                                                                      --   1: Enable Circulate  when 1;     0: send fifo data only once
                                                                      --   2: Enable Triggered Mode when 1; 0: run continueously (no TTC)
                                                                      --   3: Enable pattern generator
                                                                      
  end record;

  type bitfield_mrod_tcvrctrl_w_type is record
    SLIDEMAX                       : std_logic_vector(23 downto 16);  -- Maximum RXSLIDES before fire a TCVR reset
    SLIDEWAIT                      : std_logic_vector(15 downto 8);   -- RXclk delay in TCVR for next RX_SLIDE operation
    FRAMESIZE                      : std_logic_vector(7 downto 0);    -- Number of 32 data words in 1 frame
  end record;


  -- Control Record
  type register_map_control_type is record
    STATUS_LEDS                    : std_logic_vector(7 downto 0);    -- Board GPIO Leds
    TIMEOUT_CTRL                   : bitfield_timeout_ctrl_w_type;   -- Central Router ToHost Controls and Monitors 
    CRTOHOST_FIFO_STATUS           : bitfield_crtohost_fifo_status_t_type;  -- Central Router ToHost Controls and Monitors 
    CRTOHOST_DMA_DESCRIPTOR_1      : bitfield_crtohost_dma_descriptor_1_t_type;  -- Central Router ToHost Controls and Monitors 
    CRTOHOST_DMA_DESCRIPTOR_2      : bitfield_crtohost_dma_descriptor_2_w_type;  -- Central Router ToHost Controls and Monitors 
    CRFROMHOST_FIFO_STATUS         : bitfield_crfromhost_fifo_status_t_type;  -- Central Router FromHost Controls and Monitors 
    BROADCAST_ENABLE               : bitfield_broadcast_enable_w_array_type; -- Enable path to be included in a broadcast message.
    CRFROMHOST_RESET               : std_logic_vector(64 downto 64);  -- Central Router FromHost Controls and Monitors
    HAS_STREAM_ID                  : bitfield_has_stream_id_w_array_type; -- Decoding block
    DECODING_EGROUP_CTRL           : bitfield_decoding_egroup_ctrl_w_2d_array_type;  -- Contols Egroup for lpGBT and GBT based links 
    MINI_EGROUP_TOHOST             : bitfield_mini_egroup_tohost_w_array_type; -- Configures the ToHost Mini egroup
    TTC_TOHOST_ENABLE              : std_logic_vector(0 downto 0);    -- Enables the ToHost Mini Egroup in TTC mode
    DECODING_REVERSE_10B           : std_logic_vector(0 downto 0);    -- Reverse 10-bit word of elink data for 8b10b E-links
                                                                      -- 1: Receive 10-bit word in ToHost E-Paths, MSB first
                                                                      -- 0: Receive 10-bit word in ToHost E-Paths, LSB first
                                                                      
    YARR_DEBUG_ALLEGROUP_TOHOST    : bitfield_yarr_debug_allegroup_tohost_w_array_type; -- Decoding block
    SUPER_CHUNK_FACTOR_LINK        : bitfield_super_chunk_factor_link_w_array_type; -- number of chunks glued together
    DECODING_LINK_CB               : bitfield_decoding_link_cb_w_array_type; -- Decoding block
    DECODING_MASK64B66BKBLOCK      : std_logic_vector(3 downto 0);    -- Mask User K-Block based on its block number (see sp011)
    DECODING_DISEGROUP             : std_logic_vector(6 downto 0);    -- Disable egroups for debugging purposes
    FULLMODE_32B_SOP               : std_logic_vector(0 downto 0);    -- When set to 1, use 32-bit 0x0000003C as start of chunk, otherwise only 8-bit 0x3C (FULL mode only)
    ENCODING_REVERSE_10B           : std_logic_vector(0 downto 0);    -- Reverse 10-bit word of elink data for 8b10b E-links. 1 MSB first, 0 LSB first
    ENCODING_EGROUP_CTRL           : bitfield_encoding_egroup_ctrl_w_2d_array_type;  -- See Central Router Doc, indices [3,4] are optimized out in wideMode 
    MINI_EGROUP_FROMHOST           : bitfield_mini_egroup_fromhost_w_array_type; -- Configures the FromHost Mini egroup
    ENCODING_EGROUP_FEI4_CTRL      : bitfield_encoding_egroup_fei4_ctrl_w_2d_array_type;  -- FEI4 encoder configuration registers. 
    YARR_DEBUG_ALLEGROUP_FROMHOST1 : bitfield_yarr_debug_allegroup_fromhost1_w_array_type; -- Encoding block
    YARR_DEBUG_ALLEGROUP_FROMHOST2 : bitfield_yarr_debug_allegroup_fromhost2_w_array_type; -- Encoding block
    YARR_FROMHOST_CALTRIGSEQ_WE    : std_logic_vector(0 downto 0);    -- enable to store CalPulse+Trigger Sequence into memory
    YARR_FROMHOST_CALTRIGSEQ_WRDATA : std_logic_vector(15 downto 0);   -- CalPulse+Trigger Sequence to be stored in memory
    YARR_FROMHOST_CALTRIGSEQ_WRADDR : std_logic_vector(4 downto 0);    -- memory address to store CalPulse+Trigger Sequence
    FE_EMU_ENA                     : bitfield_fe_emu_ena_w_type;     -- Frontend Emulator Controls and Monitors 
    FE_EMU_CONFIG                  : bitfield_fe_emu_config_w_type;  -- Frontend Emulator Controls and Monitors 
    FE_EMU_READ                    : bitfield_fe_emu_read_w_type;    -- Frontend Emulator Controls and Monitors 
    FE_EMU_LOGIC                   : bitfield_fe_emu_logic_w_type;   -- Frontend Emulator Controls and Monitors 
    GBT_CHANNEL_DISABLE            : std_logic_vector(47 downto 0);   -- Disable selected lpGBT, GBT or FULL mode channel
    GBT_GENERAL_CTRL               : std_logic_vector(63 downto 0);   -- Alignment chk reset (not self clearing)
    GBT_MODE_CTRL                  : bitfield_gbt_mode_ctrl_w_type;  -- Link Wrapper Controls 
    GBT_RXSLIDE_SELECT             : std_logic_vector(47 downto 0);   -- RxSlide select [47:0]
    GBT_RXSLIDE_MANUAL             : std_logic_vector(47 downto 0);   -- RxSlide select [47:0]
    GBT_TXUSRRDY                   : std_logic_vector(47 downto 0);   -- TxUsrRdy [47:0]
    GBT_RXUSRRDY                   : std_logic_vector(47 downto 0);   -- RxUsrRdy [47:0]
    GBT_SOFT_RESET                 : std_logic_vector(47 downto 0);   -- SOFT_RESET [47:0]
    GBT_GTTX_RESET                 : std_logic_vector(47 downto 0);   -- GTTX_RESET [47:0]
    GBT_GTRX_RESET                 : std_logic_vector(47 downto 0);   -- GTRX_RESET [47:0]
    GBT_PLL_RESET                  : bitfield_gbt_pll_reset_w_type;  -- Link Wrapper Controls 
    GBT_SOFT_TX_RESET              : bitfield_gbt_soft_tx_reset_w_type;  -- Link Wrapper Controls 
    GBT_SOFT_RX_RESET              : bitfield_gbt_soft_rx_reset_w_type;  -- Link Wrapper Controls 
    GBT_ODD_EVEN                   : std_logic_vector(47 downto 0);   -- OddEven [47:0]
    GBT_TOPBOT                     : std_logic_vector(47 downto 0);   -- TopBot [47:0]
    GBT_TX_TC_DLY_VALUE1           : std_logic_vector(47 downto 0);   -- TX_TC_DLY_VALUE [47:0]
    GBT_TX_TC_DLY_VALUE2           : std_logic_vector(47 downto 0);   -- TX_TC_DLY_VALUE [95:48]
    GBT_TX_TC_DLY_VALUE3           : std_logic_vector(47 downto 0);   -- TX_TC_DLY_VALUE [143:96]
    GBT_TX_TC_DLY_VALUE4           : std_logic_vector(47 downto 0);   -- TX_TC_DLY_VALUE [191:144]
    GBT_DATA_TXFORMAT1             : std_logic_vector(47 downto 0);   -- DATA_TXFORMAT [47:0]
    GBT_DATA_TXFORMAT2             : std_logic_vector(47 downto 0);   -- DATA_TXFORMAT [95:48]
    GBT_DATA_RXFORMAT1             : std_logic_vector(47 downto 0);   -- DATA_RXFORMAT [47:0]
    GBT_DATA_RXFORMAT2             : std_logic_vector(47 downto 0);   -- DATA_RXFORMAT [95:0]
    GBT_TX_RESET                   : std_logic_vector(47 downto 0);   -- TX Logic reset [47:0]
    GBT_RX_RESET                   : std_logic_vector(47 downto 0);   -- RX Logic reset [47:0]
    GBT_TX_TC_METHOD               : std_logic_vector(47 downto 0);   -- TX time domain crossing method [47:0]
    GBT_OUTMUX_SEL                 : std_logic_vector(47 downto 0);   -- Descrambler output MUX selection [47:0]
    GBT_TC_EDGE                    : std_logic_vector(47 downto 0);   -- Sampling edge selection for TX domain crossing [47:0]
    GBT_TXPOLARITY                 : std_logic_vector(47 downto 0);   -- 0: default polarity
                                                                      -- 1: reversed polarity for transmitter of GTH channels
                                                                      
    GBT_RXPOLARITY                 : std_logic_vector(47 downto 0);   -- 0: default polarity
                                                                      -- 1: reversed polarity for the receiver of the GTH channels
                                                                      
    GTH_LOOPBACK_CONTROL           : std_logic_vector(2 downto 0);    -- Controls loopback  for loopback: read UG476 for the details. NOTE: the TXBUFFER is disabled, near end PCS loopback is not supported.
                                                                      --   000: Normal operation
                                                                      --   001: Near-End PCS Loopback
                                                                      --   010: Near-End PMA Loopback
                                                                      --   011: Reserved
                                                                      --   100: Far-End PMA Loopback
                                                                      --   101: Reserved
                                                                      --   110: Far-End PCS Loopback 
                                                                      
    LPGBT_FEC                      : std_logic_vector(47 downto 0);   -- 0: FEC5 
                                                                      -- 1: FEC12
                                                                      
    LPGBT_DATARATE                 : std_logic_vector(47 downto 0);   -- 0: 10.24 Gbps 
                                                                      -- 1: 5.12 Gbps
                                                                      
    GBT_TOHOST_FANOUT              : bitfield_gbt_tohost_fanout_w_type;  -- Link Wrapper Controls 
    GBT_TOFRONTEND_FANOUT          : bitfield_gbt_tofrontend_fanout_w_type;  -- Link Wrapper Controls 
    FULLMODE_AUTO_RX_RESET         : bitfield_fullmode_auto_rx_reset_w_type;  -- Link Wrapper Controls 
    TTC_DEC_CTRL                   : bitfield_ttc_dec_ctrl_w_type;   -- TTC and BUSY Controls and Monitors 
    TTC_EMU                        : bitfield_ttc_emu_w_type;        -- TTC and BUSY Controls and Monitors 
    TTC_DELAY                      : std_logic_vector(3 downto 0);    -- Controls the TTC Fanout delay value, in 25ns (1BC) units
    TTC_BUSY_TIMING_CTRL           : bitfield_ttc_busy_timing_ctrl_w_type;  -- TTC and BUSY Controls and Monitors 
    TTC_BUSY_CLEAR                 : std_logic_vector(64 downto 64);  -- clears the latching busy bits in TTC_BUSY_ACCEPTED
    TTC_EMU_CONTROL                : bitfield_ttc_emu_control_w_type;  -- TTC and BUSY Controls and Monitors 
    TTC_EMU_L1A_PERIOD             : std_logic_vector(31 downto 0);   -- L1A period in BC. 0 means manual L1A with TTC_EMU_CONTROL.L1A
    TTC_EMU_ECR_PERIOD             : std_logic_vector(31 downto 0);   -- ECR period in BC. 0 means manual ECR with TTC_EMU_CONTROL.ECR
    TTC_EMU_BCR_PERIOD             : std_logic_vector(31 downto 0);   -- BCR period in BC. 0 means manual BCR with TTC_EMU_CONTROL.BCR
    TTC_EMU_LONG_CHANNEL_DATA      : std_logic_vector(31 downto 0);   -- Long channel data for the TTC emulator
    TTC_EMU_RESET                  : std_logic_vector(64 downto 64);  -- Any write to this register resets the TTC Emulator to the default state.
    TTC_ECR_MONITOR                : bitfield_ttc_ecr_monitor_t_type;  -- Counts the number of ECRs received from the TTC system, any write to this register clears the counter 
    TTC_TTYPE_MONITOR              : bitfield_ttc_ttype_monitor_t_type;  -- Counts the number of TType received from the TTC system, any write to this register clears the counter 
    TTC_BCR_PERIODICITY_MONITOR    : bitfield_ttc_bcr_periodicity_monitor_t_type;  -- Counts the number of times the BCR period does not match 3564, any write to this register clears the counter 
    TTC_BCR_COUNTER                : bitfield_ttc_bcr_counter_t_type;  -- Counts the number of times BCR is issued, any write to this register clears the counter 
    XOFF_FM_CH_FIFO_THRESH_LOW     : std_logic_vector(3 downto 0);    -- Controls the low threshold of the channel fifo in FULL mode on which
                                                                      -- an Xon will be asserted, bitfields control 4 MSB
                                                                      
    XOFF_FM_CH_FIFO_THRESH_HIGH    : std_logic_vector(3 downto 0);    -- Controls the high threshold of the channel fifo in FULL mode on which
                                                                      -- an Xoff will be asserted, bitfields control 4 MSB
                                                                      
    XOFF_FM_HIGH_THRESH            : bitfield_xoff_fm_high_thresh_t_type;  -- XOFF Controls and Monitors, see table 2 of Busy specs manual 
    XOFF_FM_SOFT_XOFF              : std_logic_vector(23 downto 0);   -- Set any bit in this register to assert XOFF for the given channel, clearing bits will assert XON
    XOFF_ENABLE                    : std_logic_vector(23 downto 0);   -- Enable XOFF assertion (To Frontend) in case the FULL mode CH FIFO gets beyond thresholds. One bit per channel
    DMA_BUSY_STATUS                : bitfield_dma_busy_status_t_type;  -- XOFF Controls and Monitors, see table 2 of Busy specs manual 
    FM_BUSY_CHANNEL_STATUS         : bitfield_fm_busy_channel_status_t_type;  -- XOFF Controls and Monitors, see table 2 of Busy specs manual 
    BUSY_MAIN_OUTPUT_FIFO_THRESH   : bitfield_busy_main_output_fifo_thresh_w_type;  -- XOFF Controls and Monitors, see table 2 of Busy specs manual 
    BUSY_MAIN_OUTPUT_FIFO_STATUS   : bitfield_busy_main_output_fifo_status_t_type;  -- XOFF Controls and Monitors, see table 2 of Busy specs manual 
    ELINK_BUSY_ENABLE              : bitfield_elink_busy_enable_w_array_type; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
    BUSY_TOHOST_ENABLE             : std_logic_vector(0 downto 0);    -- Enable the busy ToHost Virtual Elink
    HK_CTRL_I2C                    : bitfield_hk_ctrl_i2c_w_type;    -- House Keeping Controls and Monitors 
    HK_CTRL_FMC                    : bitfield_hk_ctrl_fmc_w_type;    -- House Keeping Controls and Monitors 
    HK_MON_FMC                     : bitfield_hk_mon_fmc_w_type;     -- House Keeping Controls and Monitors 
    MMCM_MAIN                      : bitfield_mmcm_main_w_type;      -- House Keeping Controls and Monitors 
    I2C_WR                         : bitfield_i2c_wr_t_type;         -- House Keeping Controls and Monitors 
    I2C_RD                         : bitfield_i2c_rd_t_type;         -- House Keeping Controls and Monitors 
    INT_TEST                       : bitfield_int_test_t_type;       -- House Keeping Controls and Monitors 
    CONFIG_FLASH_WR                : bitfield_config_flash_wr_w_type;  -- House Keeping Controls and Monitors 
    RXUSRCLK_FREQ                  : bitfield_rxusrclk_freq_w_type;  -- House Keeping Controls and Monitors 
    FELIG_L1ID_RESET               : std_logic_vector(64 downto 64);  -- Any write to this register clears the FELIG L1ID
    FELIG_DATA_GEN_CONFIG          : bitfield_felig_data_gen_config_w_array_type; -- FELIG specific configuration test registers
    FELIG_ELINK_CONFIG             : bitfield_felig_elink_config_w_array_type; -- FELIG specific configuration test registers
    FELIG_ELINK_ENABLE             : bitfield_felig_elink_enable_w_array_type; -- FELIG specific configuration registers
    FELIG_GLOBAL_CONTROL           : bitfield_felig_global_control_w_type;  -- Specific registers for Hardware based Generators 
    FELIG_LANE_CONFIG              : bitfield_felig_lane_config_w_array_type; -- FELIG specific configuration registers
    FELIG_MON_FREQ_GLOBAL          : bitfield_felig_mon_freq_global_w_type;  -- Specific registers for Hardware based Generators 
    FELIG_RESET                    : bitfield_felig_reset_w_type;    -- Specific registers for Hardware based Generators 
    FELIG_RX_SLIDE_RESET           : std_logic_vector(23 downto 0);   -- One bit per lane.  When set to 1, resets the gbt rx slide counter.
    FELIG_ITK_STRIPS_DATA_GEN_CONFIG : bitfield_felig_itk_strips_data_gen_config_w_array_type; -- ITk Strips emulator specific configuration test registers
    FMEMU_COUNTERS                 : bitfield_fmemu_counters_w_type;  -- Specific registers for Hardware based Generators 
    FMEMU_CONTROL                  : bitfield_fmemu_control_w_type;  -- Specific registers for Hardware based Generators 
    FMEMU_RANDOM_RAM_ADDR          : std_logic_vector(9 downto 0);    -- Controls the address of the ramblock for the random number generator
    FMEMU_RANDOM_RAM               : bitfield_fmemu_random_ram_t_type;  -- Specific registers for Hardware based Generators 
    FMEMU_RANDOM_CONTROL           : bitfield_fmemu_random_control_w_type;  -- Controls the random chunk length generator 
    FMEMU_CONFIG_WRADDR            : std_logic_vector(9 downto 0);    -- write enable for the FMEmu ram block
    FMEMU_CONFIG                   : bitfield_fmemu_config_t_type;   -- Specific registers for Hardware based Generators 
    WISHBONE_CONTROL               : bitfield_wishbone_control_w_type;  -- Wishbone 
    WISHBONE_WRITE                 : bitfield_wishbone_write_t_type;  -- Wishbone 
    WISHBONE_READ                  : bitfield_wishbone_read_t_type;  -- Wishbone 
    IPBUS_WRITE_ADDRESS            : std_logic_vector(31 downto 0);   -- Address of the IPBus Write RAM
    IPBUS_WRITE_DATA               : bitfield_ipbus_write_data_t_type;  -- IPbus data to write to RAM 
    IPBUS_READ_ADDRESS             : std_logic_vector(31 downto 0);   -- Address of the IPBus Read RAM
    GLOBAL_STRIPS_CONFIG           : bitfield_global_strips_config_w_type;  -- Configuration affecting all Strips links on this FELIX device 
    GLOBAL_TRICKLE_TRIGGER         : std_logic_vector(64 downto 64);  -- writing to this register issues a single trickle trigger for every LCB link connected to this FELIX device
    STRIPS_R3_TRIGGER              : std_logic_vector(64 downto 64);  -- (for tests only) simulate R3 trigger (issues 4-5 sequential triggers)
    STRIPS_L1_TRIGGER              : std_logic_vector(64 downto 64);  -- (for tests only) simulate L1 trigger (issues 4-5 sequential triggers)
    STRIPS_R3L1_TRIGGER            : std_logic_vector(64 downto 64);  -- (for tests only) simulate simultaneous R3 and L1 trigger (issues 4-5 sequential triggers)
    MROD_CTRL                      : bitfield_mrod_ctrl_w_type;      -- Specific registers for MROD 
    MROD_TCVRCTRL                  : bitfield_mrod_tcvrctrl_w_type;  -- Specific registers for MROD 
    MROD_EP0_CSMENABLE             : std_logic_vector(23 downto 0);   -- EP0 CSM Data Enable channel 23-0
    MROD_EP0_EMPTYSUPPR            : std_logic_vector(23 downto 0);   -- EP0 Set Empty Suppression channel 23-0
    MROD_EP0_HPTDCMODE             : std_logic_vector(23 downto 0);   -- EP0 Set HPTDC Mode channel 23-0
    MROD_EP0_CLRFIFOS              : std_logic_vector(23 downto 0);   -- EP0 Clear FIFOs channel 23-0
    MROD_EP0_EMULOADENA            : std_logic_vector(23 downto 0);   -- EP0 Emulator Load Enable channel 23-0
    MROD_EP0_TRXLOOPBACK           : std_logic_vector(23 downto 0);   -- EP0 Transceiver Loopback Enable channel 23-0
    MROD_EP0_TXCVRRESET            : std_logic_vector(23 downto 0);   -- EP0 Transceiver Reset all channel 23-0
    MROD_EP0_RXRESET               : std_logic_vector(23 downto 0);   -- EP0 Receiver Reset channel 23-0
    MROD_EP0_TXRESET               : std_logic_vector(23 downto 0);   -- EP0 Transmitter Reset channel 23-0
    MROD_EP1_CSMENABLE             : std_logic_vector(23 downto 0);   -- EP1 CSM Data Enable channel 23-0
    MROD_EP1_EMPTYSUPPR            : std_logic_vector(23 downto 0);   -- EP1 Set Empty Suppression channel 23-0
    MROD_EP1_HPTDCMODE             : std_logic_vector(23 downto 0);   -- EP1 Set HPTDC Mode channel 23-0
    MROD_EP1_CLRFIFOS              : std_logic_vector(23 downto 0);   -- EP1 Clear FIFOs channel 23-0
    MROD_EP1_EMULOADENA            : std_logic_vector(23 downto 0);   -- EP1 Emulator Load Enable channel 23-0
    MROD_EP1_TRXLOOPBACK           : std_logic_vector(23 downto 0);   -- EP1 Transceiver Loopback Enable channel 23-0
    MROD_EP1_TXCVRRESET            : std_logic_vector(23 downto 0);   -- EP1 Transceiver Reset all channel 23-0
    MROD_EP1_RXRESET               : std_logic_vector(23 downto 0);   -- EP1 Receiver Reset channel 23-0
    MROD_EP1_TXRESET               : std_logic_vector(23 downto 0);   -- EP1 Transmitter Reset channel 23-0
  end record;
  -----------------------------------
  ---- GENERATED code END #2 ##  ----
  -----------------------------------

  constant REG_BUSY_THRESH_ASSERT_C : std_logic_vector(63 downto 0) := x"0000_0000_0C80_0000"; --200 MB busy threshold default value.
  constant REG_BUSY_THRESH_NEGATE_C : std_logic_vector(63 downto 0) := x"0000_0000_0DC0_0000"; --220 MB busy threshold default value.

  --!
  --! --> Read/Write User Application Registers DEFAULT values (Written by PCIe)
  ------------------------------------
  ---- ## GENERATED code BEGIN #3 ----
  ------------------------------------
  constant REG_STATUS_LEDS_C                       : std_logic_vector(7 downto 0)     := x"ab";                 -- Board GPIO Leds
  constant REG_TIMEOUT_CTRL_ENABLE_C               : std_logic_vector(32 downto 32)   := "1";                   -- 1 enables the timout trailer generation for ToHost mode
  constant REG_TIMEOUT_CTRL_TIMEOUT_C              : std_logic_vector(31 downto 0)    := x"ffffffff";           -- Number of 40 MHz clock cycles after which a timeout occurs.
  constant REG_CRTOHOST_FIFO_STATUS_CLEAR_C        : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register clears the latched FULL flags
  constant REG_CRTOHOST_DMA_DESCRIPTOR_1_WR_EN_C   : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register assigns the DMA ID to the AXIS_ID set in CRTOHOST_DMA_DESCRIPTOR_2.AXIS_ID
  constant REG_CRTOHOST_DMA_DESCRIPTOR_1_DESCR_C   : std_logic_vector(2 downto 0)     := "000";                 -- Target descriptor
  constant REG_CRTOHOST_DMA_DESCRIPTOR_2_AXIS_ID_C : std_logic_vector(10 downto 0)    := "00000000000";         -- ID of the AXI stream (E-Path ID) to associate with CRTOHOST_DMA_DESCRIPTOR_1.DESCR
  constant REG_CRFROMHOST_FIFO_STATUS_CLEAR_C      : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register clears the latched FULL flags
  constant REG_BROADCAST_ENABLE_00_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_01_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_02_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_03_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_04_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_05_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_06_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_07_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_08_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_09_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_10_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_11_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_12_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_13_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_14_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_15_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_16_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_17_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_18_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_19_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_20_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_21_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_22_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_BROADCAST_ENABLE_23_C               : std_logic_vector(41 downto 0)    := "000000000000000000000000000000000000000000"; -- Enable path to be included in a broadcast message.
  constant REG_CRFROMHOST_RESET_C                  : std_logic_vector(64 downto 64)   := "0";                   -- Central Router FromHost Controls and Monitors
  constant REG_LINK_00_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_00_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_00_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_00_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_00_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_00_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_00_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_01_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_01_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_01_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_01_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_01_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_01_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_01_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_02_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_02_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_02_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_02_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_02_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_02_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_02_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_03_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_03_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_03_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_03_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_03_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_03_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_03_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_04_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_04_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_04_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_04_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_04_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_04_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_04_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_05_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_05_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_05_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_05_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_05_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_05_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_05_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_06_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_06_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_06_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_06_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_06_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_06_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_06_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_07_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_07_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_07_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_07_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_07_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_07_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_07_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_08_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_08_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_08_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_08_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_08_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_08_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_08_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_09_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_09_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_09_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_09_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_09_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_09_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_09_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_10_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_10_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_10_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_10_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_10_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_10_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_10_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_11_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_11_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_11_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_11_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_11_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_11_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_11_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_12_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_12_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_12_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_12_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_12_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_12_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_12_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_13_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_13_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_13_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_13_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_13_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_13_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_13_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_14_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_14_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_14_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_14_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_14_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_14_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_14_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_15_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_15_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_15_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_15_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_15_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_15_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_15_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_16_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_16_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_16_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_16_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_16_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_16_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_16_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_17_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_17_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_17_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_17_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_17_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_17_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_17_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_18_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_18_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_18_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_18_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_18_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_18_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_18_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_19_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_19_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_19_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_19_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_19_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_19_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_19_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_20_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_20_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_20_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_20_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_20_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_20_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_20_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_21_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_21_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_21_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_21_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_21_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_21_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_21_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_22_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_22_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_22_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_22_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_22_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_22_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_22_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_LINK_23_HAS_STREAM_ID_EGROUP6_C     : std_logic_vector(55 downto 48)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_23_HAS_STREAM_ID_EGROUP5_C     : std_logic_vector(47 downto 40)   := x"00";                 -- EPATH (Wide mode or lpGBT) is associated with a STREAM ID
  constant REG_LINK_23_HAS_STREAM_ID_EGROUP4_C     : std_logic_vector(39 downto 32)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_23_HAS_STREAM_ID_EGROUP3_C     : std_logic_vector(31 downto 24)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_23_HAS_STREAM_ID_EGROUP2_C     : std_logic_vector(23 downto 16)   := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_23_HAS_STREAM_ID_EGROUP1_C     : std_logic_vector(15 downto 8)    := x"00";                 -- EPATH is associated with a STREAM ID
  constant REG_LINK_23_HAS_STREAM_ID_EGROUP0_C     : std_logic_vector(7 downto 0)     := x"00";                 -- EPATH is associated with a STREAM ID, use only bit0 for FULL mode.
  constant REG_DECODING_LINK00_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK00_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK00_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK00_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK00_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK00_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK00_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK00_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK00_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK00_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK00_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK00_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK00_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK00_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK00_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK00_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK00_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK00_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK00_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK00_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK00_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK00_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK00_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK00_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK00_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK00_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK00_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK00_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK00_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK00_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK00_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK00_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK00_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK00_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK00_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK01_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK01_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK01_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK01_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK01_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK01_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK01_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK01_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK01_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK01_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK01_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK01_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK01_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK01_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK01_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK01_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK01_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK01_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK01_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK01_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK01_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK01_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK01_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK01_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK01_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK01_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK01_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK01_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK01_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK01_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK01_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK01_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK01_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK01_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK01_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK02_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK02_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK02_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK02_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK02_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK02_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK02_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK02_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK02_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK02_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK02_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK02_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK02_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK02_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK02_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK02_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK02_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK02_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK02_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK02_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK02_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK02_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK02_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK02_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK02_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK02_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK02_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK02_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK02_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK02_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK02_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK02_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK02_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK02_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK02_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK03_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK03_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK03_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK03_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK03_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK03_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK03_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK03_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK03_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK03_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK03_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK03_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK03_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK03_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK03_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK03_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK03_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK03_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK03_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK03_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK03_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK03_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK03_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK03_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK03_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK03_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK03_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK03_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK03_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK03_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK03_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK03_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK03_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK03_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK03_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK04_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK04_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK04_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK04_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK04_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK04_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK04_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK04_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK04_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK04_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK04_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK04_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK04_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK04_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK04_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK04_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK04_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK04_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK04_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK04_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK04_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK04_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK04_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK04_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK04_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK04_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK04_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK04_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK04_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK04_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK04_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK04_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK04_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK04_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK04_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK05_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK05_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK05_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK05_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK05_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK05_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK05_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK05_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK05_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK05_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK05_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK05_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK05_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK05_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK05_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK05_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK05_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK05_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK05_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK05_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK05_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK05_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK05_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK05_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK05_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK05_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK05_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK05_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK05_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK05_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK05_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK05_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK05_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK05_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK05_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK06_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK06_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK06_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK06_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK06_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK06_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK06_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK06_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK06_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK06_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK06_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK06_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK06_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK06_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK06_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK06_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK06_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK06_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK06_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK06_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK06_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK06_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK06_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK06_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK06_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK06_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK06_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK06_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK06_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK06_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK06_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK06_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK06_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK06_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK06_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK07_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK07_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK07_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK07_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK07_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK07_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK07_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK07_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK07_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK07_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK07_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK07_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK07_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK07_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK07_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK07_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK07_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK07_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK07_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK07_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK07_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK07_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK07_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK07_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK07_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK07_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK07_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK07_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK07_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK07_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK07_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK07_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK07_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK07_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK07_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK08_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK08_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK08_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK08_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK08_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK08_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK08_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK08_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK08_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK08_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK08_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK08_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK08_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK08_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK08_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK08_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK08_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK08_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK08_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK08_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK08_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK08_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK08_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK08_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK08_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK08_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK08_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK08_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK08_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK08_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK08_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK08_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK08_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK08_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK08_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK09_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK09_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK09_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK09_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK09_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK09_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK09_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK09_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK09_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK09_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK09_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK09_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK09_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK09_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK09_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK09_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK09_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK09_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK09_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK09_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK09_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK09_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK09_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK09_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK09_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK09_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK09_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK09_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK09_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK09_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK09_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK09_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK09_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK09_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK09_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK10_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK10_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK10_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK10_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK10_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK10_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK10_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK10_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK10_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK10_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK10_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK10_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK10_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK10_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK10_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK10_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK10_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK10_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK10_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK10_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK10_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK10_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK10_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK10_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK10_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK10_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK10_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK10_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK10_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK10_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK10_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK10_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK10_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK10_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK10_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK11_EGROUP0_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK11_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK11_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK11_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK11_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK11_EGROUP1_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK11_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK11_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK11_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK11_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK11_EGROUP2_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK11_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK11_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK11_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK11_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK11_EGROUP3_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK11_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK11_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK11_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK11_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK11_EGROUP4_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK11_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK11_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK11_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK11_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK11_EGROUP5_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK11_EGROUP5_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK11_EGROUP5_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK11_EGROUP5_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK11_EGROUP5_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_DECODING_LINK11_EGROUP6_CTRL_ENABLE_TRUNCATION_C: std_logic_vector(59 downto 59)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_DECODING_LINK11_EGROUP6_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_DECODING_LINK11_EGROUP6_CTRL_PATH_ENCODING_C: std_logic_vector(42 downto 11)   := x"11111111";           -- Encoding for every EPATH, 4 bits per E-path
                                                                                                                -- 0: direct mode
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: TTC
                                                                                                                -- 4: ITk Strips 8b10b
                                                                                                                -- 5: ITk Pixel
                                                                                                                -- 6: Endeavour
                                                                                                                -- 7-15:  reserved
                                                                                                                
  constant REG_DECODING_LINK11_EGROUP6_CTRL_EPATH_WIDTH_C: std_logic_vector(10 downto 8)    := "000";                 -- Width in bits of all EPATHS in an EGROUP 0:2, 1:4, 2:8, 3:16, 4:32
  constant REG_DECODING_LINK11_EGROUP6_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per EPATH
  constant REG_MINI_EGROUP_TOHOST_00_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_00_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_00_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_00_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_00_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_00_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_00_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_00_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_00_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_00_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_01_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_01_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_01_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_01_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_01_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_01_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_01_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_01_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_01_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_01_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_02_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_02_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_02_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_02_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_02_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_02_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_02_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_02_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_02_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_02_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_03_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_03_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_03_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_03_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_03_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_03_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_03_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_03_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_03_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_03_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_04_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_04_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_04_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_04_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_04_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_04_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_04_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_04_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_04_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_04_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_05_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_05_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_05_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_05_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_05_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_05_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_05_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_05_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_05_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_05_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_06_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_06_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_06_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_06_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_06_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_06_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_06_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_06_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_06_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_06_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_07_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_07_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_07_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_07_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_07_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_07_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_07_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_07_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_07_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_07_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_08_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_08_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_08_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_08_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_08_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_08_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_08_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_08_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_08_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_08_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_09_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_09_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_09_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_09_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_09_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_09_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_09_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_09_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_09_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_09_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_10_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_10_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_10_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_10_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_10_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_10_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_10_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_10_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_10_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_10_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_11_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_11_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_11_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_11_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_11_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_11_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_11_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_11_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_11_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_11_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_12_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_12_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_12_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_12_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_12_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_12_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_12_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_12_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_12_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_12_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_13_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_13_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_13_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_13_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_13_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_13_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_13_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_13_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_13_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_13_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_14_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_14_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_14_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_14_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_14_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_14_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_14_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_14_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_14_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_14_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_15_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_15_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_15_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_15_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_15_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_15_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_15_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_15_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_15_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_15_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_16_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_16_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_16_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_16_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_16_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_16_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_16_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_16_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_16_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_16_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_17_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_17_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_17_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_17_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_17_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_17_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_17_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_17_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_17_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_17_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_18_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_18_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_18_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_18_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_18_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_18_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_18_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_18_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_18_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_18_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_19_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_19_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_19_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_19_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_19_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_19_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_19_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_19_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_19_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_19_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_20_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_20_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_20_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_20_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_20_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_20_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_20_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_20_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_20_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_20_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_21_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_21_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_21_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_21_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_21_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_21_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_21_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_21_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_21_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_21_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_22_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_22_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_22_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_22_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_22_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_22_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_22_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_22_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_22_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_22_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_MINI_EGROUP_TOHOST_23_ENABLE_AUX_TRUNCATION_C: std_logic_vector(15 downto 15)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_23_ENABLE_IC_TRUNCATION_C: std_logic_vector(14 downto 14)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_23_ENABLE_EC_TRUNCATION_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable truncation mechanism in HDLC decoder for chunks > 12 bytes
  constant REG_MINI_EGROUP_TOHOST_23_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_23_AUX_ENABLE_C  : std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_TOHOST_23_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_23_IC_ENABLE_C   : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_TOHOST_23_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two input bits of EC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_TOHOST_23_EC_ENCODING_C : std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_TOHOST_23_EC_ENABLE_C   : std_logic_vector(0 downto 0)     := "1";                   -- Enables the EC channel
  constant REG_TTC_TOHOST_ENABLE_C                 : std_logic_vector(0 downto 0)     := "1";                   -- Enables the ToHost Mini Egroup in TTC mode
  constant REG_DECODING_REVERSE_10B_C              : std_logic_vector(0 downto 0)     := "1";                   -- Reverse 10-bit word of elink data for 8b10b E-links
                                                                                                                -- 1: Receive 10-bit word in ToHost E-Paths, MSB first
                                                                                                                -- 0: Receive 10-bit word in ToHost E-Paths, LSB first
                                                                                                                
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_00_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_01_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_02_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_03_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_04_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_05_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_06_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_07_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_08_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_09_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_10_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_YARR_DEBUG_ALLEGROUP_TOHOST_11_REF_PACKET_C: std_logic_vector(63 downto 32)   := x"02000000";           -- Reference packet to be matched
  constant REG_SUPER_CHUNK_FACTOR_LINK_00_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_01_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_02_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_03_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_04_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_05_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_06_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_07_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_08_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_09_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_10_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_SUPER_CHUNK_FACTOR_LINK_11_C        : std_logic_vector(7 downto 0)     := x"01";                 -- number of chunks glued together
  constant REG_DECODING_LINK_00_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_01_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_02_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_03_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_04_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_05_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_06_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_07_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_08_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_09_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_10_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_LINK_11_CB_CBOPT_C         : std_logic_vector(3 downto 0)     := x"0";                  -- Channel bonding option
                                                                                                                -- 0: no bonding
                                                                                                                -- 3: Bonding 0/1/2 3/4/5
                                                                                                                -- other values: reserved
                                                                                                                
  constant REG_DECODING_MASK64B66BKBLOCK_C         : std_logic_vector(3 downto 0)     := x"a";                  -- Mask User K-Block based on its block number (see sp011)
  constant REG_DECODING_DISEGROUP_C                : std_logic_vector(6 downto 0)     := "0000000";             -- Disable egroups for debugging purposes
  constant REG_FULLMODE_32B_SOP_C                  : std_logic_vector(0 downto 0)     := "0";                   -- When set to 1, use 32-bit 0x0000003C as start of chunk, otherwise only 8-bit 0x3C (FULL mode only)
  constant REG_ENCODING_REVERSE_10B_C              : std_logic_vector(0 downto 0)     := "1";                   -- Reverse 10-bit word of elink data for 8b10b E-links. 1 MSB first, 0 LSB first
  constant REG_ENCODING_LINK00_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK00_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK00_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK00_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK00_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK00_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK00_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK00_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK00_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK00_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK00_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK00_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK00_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK00_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK00_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK00_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK00_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK00_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK00_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK00_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK00_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK01_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK01_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK01_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK01_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK01_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK01_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK01_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK01_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK01_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK01_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK01_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK01_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK01_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK01_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK01_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK01_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK01_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK01_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK01_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK01_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK01_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK02_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK02_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK02_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK02_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK02_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK02_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK02_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK02_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK02_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK02_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK02_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK02_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK02_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK02_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK02_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK02_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK02_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK02_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK02_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK02_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK02_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK03_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK03_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK03_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK03_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK03_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK03_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK03_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK03_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK03_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK03_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK03_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK03_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK03_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK03_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK03_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK03_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK03_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK03_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK03_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK03_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK03_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK04_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK04_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK04_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK04_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK04_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK04_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK04_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK04_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK04_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK04_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK04_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK04_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK04_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK04_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK04_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK04_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK04_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK04_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK04_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK04_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK04_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK05_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK05_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK05_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK05_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK05_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK05_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK05_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK05_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK05_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK05_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK05_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK05_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK05_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK05_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK05_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK05_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK05_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK05_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK05_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK05_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK05_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK06_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK06_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK06_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK06_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK06_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK06_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK06_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK06_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK06_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK06_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK06_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK06_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK06_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK06_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK06_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK06_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK06_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK06_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK06_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK06_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK06_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK07_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK07_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK07_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK07_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK07_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK07_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK07_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK07_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK07_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK07_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK07_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK07_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK07_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK07_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK07_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK07_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK07_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK07_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK07_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK07_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK07_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK08_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK08_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK08_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK08_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK08_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK08_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK08_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK08_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK08_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK08_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK08_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK08_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK08_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK08_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK08_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK08_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK08_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK08_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK08_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK08_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK08_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK09_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK09_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK09_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK09_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK09_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK09_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK09_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK09_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK09_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK09_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK09_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK09_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK09_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK09_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK09_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK09_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK09_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK09_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK09_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK09_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK09_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK10_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK10_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK10_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK10_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK10_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK10_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK10_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK10_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK10_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK10_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK10_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK10_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK10_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK10_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK10_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK10_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK10_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK10_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK10_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK10_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK10_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK11_EGROUP0_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK11_EGROUP0_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK11_EGROUP0_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK11_EGROUP0_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP0_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP0_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK11_EGROUP1_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK11_EGROUP1_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK11_EGROUP1_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK11_EGROUP1_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP1_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP1_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK11_EGROUP2_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK11_EGROUP2_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK11_EGROUP2_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK11_EGROUP2_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP2_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP2_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK11_EGROUP3_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK11_EGROUP3_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK11_EGROUP3_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK11_EGROUP3_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP3_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP3_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_ENCODING_LINK11_EGROUP4_CTRL_ENABLE_DELAY_C: std_logic_vector(63 downto 63)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_ENCODING_LINK11_EGROUP4_CTRL_TTC_OPTION_C: std_logic_vector(62 downto 59)   := x"0";                  -- Selects TTC bits sent to the E-link
  constant REG_ENCODING_LINK11_EGROUP4_CTRL_REVERSE_ELINKS_C: std_logic_vector(50 downto 43)   := x"00";                 -- enables bit reversing for the elink in the given epath
  constant REG_ENCODING_LINK11_EGROUP4_CTRL_EPATH_WIDTH_C: std_logic_vector(42 downto 40)   := "000";                 -- Width of the Elinks in the egroup
                                                                                                                -- 0: 2 bit 80 Mb/s
                                                                                                                -- 1: 4 bit 160 Mb/s
                                                                                                                -- 2: 8 bit 320 Mb/s
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP4_CTRL_PATH_ENCODING_C: std_logic_vector(39 downto 8)    := x"11111111";           -- Encoding for every EPATH, 4 bits per E-Path
                                                                                                                -- 0: No encoding
                                                                                                                -- 1: 8b10b mode
                                                                                                                -- 2: HDLC mode
                                                                                                                -- 3: ITk Strip LCB
                                                                                                                -- 4: ITk Pixel
                                                                                                                -- 5: Endeavour
                                                                                                                -- 6: reserved
                                                                                                                -- 7: reserved
                                                                                                                -- greater than 7: TTC mode, see firmware Phase 2 specification doc
                                                                                                                
  constant REG_ENCODING_LINK11_EGROUP4_CTRL_EPATH_ENA_C: std_logic_vector(7 downto 0)     := x"00";                 -- Enable bits per E-PATH
  constant REG_MINI_EGROUP_FROMHOST_00_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_00_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_00_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_00_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_00_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_00_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_00_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_00_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_01_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_01_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_01_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_01_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_01_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_01_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_01_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_01_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_02_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_02_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_02_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_02_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_02_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_02_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_02_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_02_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_03_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_03_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_03_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_03_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_03_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_03_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_03_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_03_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_04_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_04_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_04_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_04_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_04_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_04_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_04_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_04_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_05_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_05_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_05_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_05_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_05_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_05_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_05_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_05_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_06_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_06_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_06_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_06_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_06_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_06_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_06_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_06_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_07_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_07_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_07_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_07_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_07_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_07_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_07_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_07_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_08_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_08_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_08_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_08_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_08_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_08_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_08_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_08_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_09_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_09_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_09_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_09_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_09_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_09_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_09_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_09_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_10_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_10_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_10_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_10_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_10_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_10_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_10_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_10_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_11_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_11_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_11_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_11_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_11_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_11_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_11_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_11_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_12_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_12_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_12_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_12_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_12_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_12_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_12_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_12_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_13_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_13_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_13_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_13_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_13_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_13_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_13_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_13_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_14_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_14_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_14_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_14_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_14_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_14_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_14_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_14_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_15_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_15_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_15_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_15_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_15_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_15_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_15_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_15_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_16_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_16_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_16_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_16_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_16_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_16_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_16_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_16_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_17_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_17_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_17_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_17_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_17_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_17_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_17_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_17_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_18_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_18_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_18_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_18_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_18_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_18_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_18_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_18_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_19_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_19_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_19_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_19_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_19_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_19_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_19_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_19_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_20_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_20_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_20_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_20_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_20_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_20_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_20_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_20_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_21_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_21_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_21_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_21_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_21_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_21_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_21_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_21_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_22_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_22_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_22_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_22_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_22_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_22_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_22_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_22_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_MINI_EGROUP_FROMHOST_23_ENABLE_DELAY_C: std_logic_vector(13 downto 13)   := "0";                   -- Enable inter-packet delay generation in HDLC encoder
  constant REG_MINI_EGROUP_FROMHOST_23_AUX_BIT_SWAPPING_C: std_logic_vector(11 downto 11)   := "1";                   -- 0: two input bits of AUX e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_23_AUX_ENABLE_C: std_logic_vector(10 downto 10)   := "1";                   -- Enables the AUX channel
  constant REG_MINI_EGROUP_FROMHOST_23_IC_BIT_SWAPPING_C: std_logic_vector(8 downto 8)     := "1";                   -- 0: two input bits of IC e-link are as documented, 1: two input bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_23_IC_ENABLE_C : std_logic_vector(7 downto 7)     := "1";                   -- Enables the IC channel
  constant REG_MINI_EGROUP_FROMHOST_23_EC_BIT_SWAPPING_C: std_logic_vector(5 downto 5)     := "0";                   -- 0: two output bits of EC e-link are as documented, 1: two output bits are swapped
  constant REG_MINI_EGROUP_FROMHOST_23_EC_ENCODING_C: std_logic_vector(4 downto 1)     := x"2";                  -- Configures encoding of the EC channel
  constant REG_MINI_EGROUP_FROMHOST_23_EC_ENABLE_C : std_logic_vector(0 downto 0)     := "1";                   -- Configures the FromHost Mini egroup
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK00_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK01_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK02_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK03_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK04_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK05_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK06_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK07_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK08_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK09_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK10_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP0_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP1_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP2_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP3_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL_PHASE_DELAY1_C: std_logic_vector(11 downto 9)    := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE1_C: std_logic_vector(8 downto 8)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE1_C: std_logic_vector(7 downto 7)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL_TTC_SELECT1_C: std_logic_vector(6 downto 6)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL_PHASE_DELAY0_C: std_logic_vector(5 downto 3)     := "000";                 -- phase delay of output data, with 320 Bb/s e-link 8 phases per BC
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL_MANCHESTER_ENABLE0_C: std_logic_vector(2 downto 2)     := "0";                   -- enable manchester encoding
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL_AUTOMATIC_MERGE_DISABLE0_C: std_logic_vector(1 downto 1)     := "0";                   -- Disable automatic merging
  constant REG_ENCODING_LINK11_EGROUP4_FEI4_CTRL_TTC_SELECT0_C: std_logic_vector(0 downto 0)     := "0";                   -- TTC/FromHost select (if automatic merging is disabled)
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_00_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_00_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_00_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_01_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_01_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_01_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_02_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_02_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_02_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_03_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_03_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_03_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_04_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_04_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_04_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_05_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_05_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_05_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_06_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_06_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_06_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_07_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_07_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_07_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_08_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_08_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_08_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_09_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_09_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_09_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_10_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_10_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_10_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_11_RD53A_AZ_EN_C: std_logic_vector(48 downto 48)   := "0";                   -- Auto zeroing module enable
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST1_11_REF_DLY_GENCALTRIG_C: std_logic_vector(7 downto 0)     := x"0f";                 -- Reference distance between GenCal and First Trigger
  constant REG_YARR_DEBUG_ALLEGROUP_FROMHOST2_11_REF_CMD_C: std_logic_vector(15 downto 0)    := x"6666";               -- Cmd type to be counted. See RD53 Manual for list of allowed commands
  constant REG_YARR_FROMHOST_CALTRIGSEQ_WE_C       : std_logic_vector(0 downto 0)     := "0";                   -- enable to store CalPulse+Trigger Sequence into memory
  constant REG_YARR_FROMHOST_CALTRIGSEQ_WRDATA_C   : std_logic_vector(15 downto 0)    := x"0000";               -- CalPulse+Trigger Sequence to be stored in memory
  constant REG_YARR_FROMHOST_CALTRIGSEQ_WRADDR_C   : std_logic_vector(4 downto 0)     := "00000";               -- memory address to store CalPulse+Trigger Sequence
  constant REG_FE_EMU_ENA_EMU_TOFRONTEND_C         : std_logic_vector(1 downto 1)     := "0";                   -- Enable GBT dummy emulator ToFrontEnd
  constant REG_FE_EMU_ENA_EMU_TOHOST_C             : std_logic_vector(0 downto 0)     := "0";                   -- Enable GBT dummy emulator ToHost
  constant REG_FE_EMU_CONFIG_WE_C                  : std_logic_vector(54 downto 47)   := x"00";                 -- write enable array, every bit is one emulator RAM block
  constant REG_FE_EMU_CONFIG_WRADDR_C              : std_logic_vector(46 downto 33)   := "00000000000000";      -- write address bus
  constant REG_FE_EMU_CONFIG_WRDATA_C              : std_logic_vector(32 downto 0)    := "000000000000000000000000000000000"; -- write data bus
  constant REG_FE_EMU_READ_SEL_C                   : std_logic_vector(35 downto 33)   := "000";                 -- Select ramblock to read back
  constant REG_FE_EMU_LOGIC_L1A_TRIGGERED_C        : std_logic_vector(33 downto 33)   := "0";                   -- 1 Send a chunk on every L1A, 0 use the IDLES to determine the rate
  constant REG_FE_EMU_LOGIC_ENA_C                  : std_logic_vector(32 downto 32)   := "0";                   -- Enable logic based FrontEnd emulator, instead of RAM based.
  constant REG_FE_EMU_LOGIC_IDLES_C                : std_logic_vector(31 downto 16)   := x"0000";               -- Number of IDLE bytes between chunks.
  constant REG_FE_EMU_LOGIC_CHUNK_LENGTH_C         : std_logic_vector(15 downto 0)    := x"0000";               -- Chunk length in bytes
  constant REG_GBT_CHANNEL_DISABLE_C               : std_logic_vector(47 downto 0)    := x"000000000000";       -- Disable selected lpGBT, GBT or FULL mode channel
  constant REG_GBT_GENERAL_CTRL_C                  : std_logic_vector(63 downto 0)    := x"0000000000000000";   -- Alignment chk reset (not self clearing)
  constant REG_GBT_MODE_CTRL_RX_ALIGN_TB_SW_C      : std_logic_vector(2 downto 2)     := "0";                   -- RX_ALIGN_TB_SW
  constant REG_GBT_MODE_CTRL_RX_ALIGN_SW_C         : std_logic_vector(1 downto 1)     := "0";                   -- RX_ALIGN_SW
  constant REG_GBT_MODE_CTRL_DESMUX_USE_SW_C       : std_logic_vector(0 downto 0)     := "0";                   -- DESMUX_USE_SW
  constant REG_GBT_RXSLIDE_SELECT_C                : std_logic_vector(47 downto 0)    := x"000000000000";       -- RxSlide select [47:0]
  constant REG_GBT_RXSLIDE_MANUAL_C                : std_logic_vector(47 downto 0)    := x"000000000000";       -- RxSlide select [47:0]
  constant REG_GBT_TXUSRRDY_C                      : std_logic_vector(47 downto 0)    := x"ffffffffffff";       -- TxUsrRdy [47:0]
  constant REG_GBT_RXUSRRDY_C                      : std_logic_vector(47 downto 0)    := x"ffffffffffff";       -- RxUsrRdy [47:0]
  constant REG_GBT_SOFT_RESET_C                    : std_logic_vector(47 downto 0)    := x"000000000000";       -- SOFT_RESET [47:0]
  constant REG_GBT_GTTX_RESET_C                    : std_logic_vector(47 downto 0)    := x"000000000000";       -- GTTX_RESET [47:0]
  constant REG_GBT_GTRX_RESET_C                    : std_logic_vector(47 downto 0)    := x"000000000000";       -- GTRX_RESET [47:0]
  constant REG_GBT_PLL_RESET_QPLL_RESET_C          : std_logic_vector(59 downto 48)   := x"000";                -- QPLL_RESET [11:0]
  constant REG_GBT_PLL_RESET_CPLL_RESET_C          : std_logic_vector(47 downto 0)    := x"000000000000";       -- CPLL_RESET [47:0]
  constant REG_GBT_SOFT_TX_RESET_RESET_ALL_C       : std_logic_vector(59 downto 48)   := x"000";                -- SOFT_TX_RESET_ALL [11:0]
  constant REG_GBT_SOFT_TX_RESET_RESET_GT_C        : std_logic_vector(47 downto 0)    := x"000000000000";       -- SOFT_TX_RESET_GT [47:0]
  constant REG_GBT_SOFT_RX_RESET_RESET_ALL_C       : std_logic_vector(59 downto 48)   := x"000";                -- SOFT_TX_RESET_ALL [11:0]
  constant REG_GBT_SOFT_RX_RESET_RESET_GT_C        : std_logic_vector(47 downto 0)    := x"000000000000";       -- SOFT_TX_RESET_GT [47:0]
  constant REG_GBT_ODD_EVEN_C                      : std_logic_vector(47 downto 0)    := x"000000000000";       -- OddEven [47:0]
  constant REG_GBT_TOPBOT_C                        : std_logic_vector(47 downto 0)    := x"000000000000";       -- TopBot [47:0]
  constant REG_GBT_TX_TC_DLY_VALUE1_C              : std_logic_vector(47 downto 0)    := x"333333333333";       -- TX_TC_DLY_VALUE [47:0]
  constant REG_GBT_TX_TC_DLY_VALUE2_C              : std_logic_vector(47 downto 0)    := x"333333333333";       -- TX_TC_DLY_VALUE [95:48]
  constant REG_GBT_TX_TC_DLY_VALUE3_C              : std_logic_vector(47 downto 0)    := x"333333333333";       -- TX_TC_DLY_VALUE [143:96]
  constant REG_GBT_TX_TC_DLY_VALUE4_C              : std_logic_vector(47 downto 0)    := x"333333333333";       -- TX_TC_DLY_VALUE [191:144]
  constant REG_GBT_DATA_TXFORMAT1_C                : std_logic_vector(47 downto 0)    := x"000000000000";       -- DATA_TXFORMAT [47:0]
  constant REG_GBT_DATA_TXFORMAT2_C                : std_logic_vector(47 downto 0)    := x"000000000000";       -- DATA_TXFORMAT [95:48]
  constant REG_GBT_DATA_RXFORMAT1_C                : std_logic_vector(47 downto 0)    := x"000000000000";       -- DATA_RXFORMAT [47:0]
  constant REG_GBT_DATA_RXFORMAT2_C                : std_logic_vector(47 downto 0)    := x"000000000000";       -- DATA_RXFORMAT [95:0]
  constant REG_GBT_TX_RESET_C                      : std_logic_vector(47 downto 0)    := x"000000000000";       -- TX Logic reset [47:0]
  constant REG_GBT_RX_RESET_C                      : std_logic_vector(47 downto 0)    := x"000000000000";       -- RX Logic reset [47:0]
  constant REG_GBT_TX_TC_METHOD_C                  : std_logic_vector(47 downto 0)    := x"000000000000";       -- TX time domain crossing method [47:0]
  constant REG_GBT_OUTMUX_SEL_C                    : std_logic_vector(47 downto 0)    := x"000000000000";       -- Descrambler output MUX selection [47:0]
  constant REG_GBT_TC_EDGE_C                       : std_logic_vector(47 downto 0)    := x"000000000000";       -- Sampling edge selection for TX domain crossing [47:0]
  constant REG_GBT_TXPOLARITY_C                    : std_logic_vector(47 downto 0)    := x"000000000000";       -- 0: default polarity
                                                                                                                -- 1: reversed polarity for transmitter of GTH channels
                                                                                                                
  constant REG_GBT_RXPOLARITY_C                    : std_logic_vector(47 downto 0)    := x"000000000000";       -- 0: default polarity
                                                                                                                -- 1: reversed polarity for the receiver of the GTH channels
                                                                                                                
  constant REG_GTH_LOOPBACK_CONTROL_C              : std_logic_vector(2 downto 0)     := "000";                 -- Controls loopback  for loopback: read UG476 for the details. NOTE: the TXBUFFER is disabled, near end PCS loopback is not supported.
                                                                                                                --   000: Normal operation
                                                                                                                --   001: Near-End PCS Loopback
                                                                                                                --   010: Near-End PMA Loopback
                                                                                                                --   011: Reserved
                                                                                                                --   100: Far-End PMA Loopback
                                                                                                                --   101: Reserved
                                                                                                                --   110: Far-End PCS Loopback 
                                                                                                                
  constant REG_LPGBT_FEC_C                         : std_logic_vector(47 downto 0)    := x"000000000000";       -- 0: FEC5 
                                                                                                                -- 1: FEC12
                                                                                                                
  constant REG_LPGBT_DATARATE_C                    : std_logic_vector(47 downto 0)    := x"000000000000";       -- 0: 10.24 Gbps 
                                                                                                                -- 1: 5.12 Gbps
                                                                                                                
  constant REG_GBT_TOHOST_FANOUT_LOCK_C            : std_logic_vector(48 downto 48)   := "0";                   -- Locks this particular register. If set prevents software from touching it.
  constant REG_GBT_TOHOST_FANOUT_SEL_C             : std_logic_vector(47 downto 0)    := x"000000000000";       -- ToHost FanOut/Selector. Every bitfield is a channel:
                                                                                                                --   1 : GBT_EMU, select GBT Emulator for a specific CentralRouter channel
                                                                                                                --   0 : GBT_WRAP, select real GBT link for a specific CentralRouter channel
                                                                                                                
  constant REG_GBT_TOFRONTEND_FANOUT_LOCK_C        : std_logic_vector(48 downto 48)   := "0";                   -- Locks this particular register. If set prevents software from touching it.
  constant REG_GBT_TOFRONTEND_FANOUT_SEL_C         : std_logic_vector(47 downto 0)    := x"000000000000";       -- ToFrontEnd FanOut/Selector. Every bitfield is a channel:
                                                                                                                --   1 : GBT_EMU, select GBT Emulator for a specific GBT link
                                                                                                                --   0 : TTC_DEC, select CentralRouter data (including TTC) for a specific GBT link
                                                                                                                --   
                                                                                                                
  constant REG_FULLMODE_AUTO_RX_RESET_ENABLE_C     : std_logic_vector(32 downto 32)   := "1";                   -- Enable the Automatic RX Reset mechanism
  constant REG_FULLMODE_AUTO_RX_RESET_TIMEOUT_C    : std_logic_vector(31 downto 0)    := x"00100000";           -- Number of 40 MHz clock cycles until an unaligned link results in a reset pulse
  constant REG_TTC_DEC_CTRL_B_CHAN_DELAY_C         : std_logic_vector(30 downto 27)   := x"0";                  -- Number of BC to delay the L1A distribution to the frontends
  constant REG_TTC_DEC_CTRL_BCID_ONBCR_C           : std_logic_vector(26 downto 15)   := x"000";                -- BCID is set to this value when BCR arrives
  constant REG_TTC_DEC_CTRL_ECR_BCR_SWAP_C         : std_logic_vector(13 downto 13)   := "0";                   -- ECR and BCR signals are swapped at the output of the TTC decoder (needed only for LAr TTC)
  constant REG_TTC_DEC_CTRL_BUSY_OUTPUT_INHIBIT_C  : std_logic_vector(12 downto 12)   := "0";                   -- forces the Busy LEMO output to BUSY-OFF
  constant REG_TTC_DEC_CTRL_TOHOST_RST_C           : std_logic_vector(11 downto 11)   := "0";                   -- reset toHost in ttc decoder
  constant REG_TTC_DEC_CTRL_TT_BCH_EN_C            : std_logic_vector(10 downto 10)   := "1";                   -- trigger type enable / disable for TTC-ToHost
  constant REG_TTC_DEC_CTRL_XL1ID_SW_C             : std_logic_vector(9 downto 2)     := x"00";                 -- set XL1ID value, the value to be set by XL1ID_RST signal
  constant REG_TTC_DEC_CTRL_XL1ID_RST_C            : std_logic_vector(1 downto 1)     := "0";                   -- giving a trigger signal to reset XL1ID value
  constant REG_TTC_DEC_CTRL_MASTER_BUSY_C          : std_logic_vector(0 downto 0)     := "0";                   -- L1A trigger throttling
  constant REG_TTC_EMU_SEL_C                       : std_logic_vector(1 downto 1)     := "0";                   -- Select TTC data source 1 TTC Emu | 0 TTC Decoder
  constant REG_TTC_EMU_ENA_C                       : std_logic_vector(0 downto 0)     := "0";                   -- Clear to load into the TTC emulator’s memory the required sequence, Set to run the TTC emulator sequence
  constant REG_TTC_DELAY_C                         : std_logic_vector(3 downto 0)     := x"0";                  -- Controls the TTC Fanout delay value, in 25ns (1BC) units
  constant REG_TTC_BUSY_TIMING_CTRL_PRESCALE_C     : std_logic_vector(51 downto 32)   := x"0000f";              -- Prescales the 40MHz clock to create an internal slow clock
  constant REG_TTC_BUSY_TIMING_CTRL_BUSY_WIDTH_C   : std_logic_vector(31 downto 16)   := x"000f";               -- Minimum number of 40MHz clocks that the busy is asserted
  constant REG_TTC_BUSY_TIMING_CTRL_LIMIT_TIME_C   : std_logic_vector(15 downto 0)    := x"000f";               -- Number of prescaled clocks a given busy must be asserted before it is recognized
  constant REG_TTC_BUSY_CLEAR_C                    : std_logic_vector(64 downto 64)   := "0";                   -- clears the latching busy bits in TTC_BUSY_ACCEPTED
  constant REG_TTC_EMU_CONTROL_BUSY_IN_ENABLE_C    : std_logic_vector(33 downto 33)   := "1";                   -- Enable internal BUSY input to stop L1A on BUSY
  constant REG_TTC_EMU_CONTROL_BROADCAST_C         : std_logic_vector(32 downto 27)   := "000000";              -- Broadcast data
  constant REG_TTC_EMU_CONTROL_ECR_C               : std_logic_vector(26 downto 26)   := "0";                   -- Event counter reset
  constant REG_TTC_EMU_CONTROL_BCR_C               : std_logic_vector(25 downto 25)   := "0";                   -- Bunch counter reset
  constant REG_TTC_EMU_CONTROL_L1A_C               : std_logic_vector(24 downto 24)   := "0";                   -- Level 1 Accept
  constant REG_TTC_EMU_L1A_PERIOD_C                : std_logic_vector(31 downto 0)    := x"00000000";           -- L1A period in BC. 0 means manual L1A with TTC_EMU_CONTROL.L1A
  constant REG_TTC_EMU_ECR_PERIOD_C                : std_logic_vector(31 downto 0)    := x"00000000";           -- ECR period in BC. 0 means manual ECR with TTC_EMU_CONTROL.ECR
  constant REG_TTC_EMU_BCR_PERIOD_C                : std_logic_vector(31 downto 0)    := x"00000dec";           -- BCR period in BC. 0 means manual BCR with TTC_EMU_CONTROL.BCR
  constant REG_TTC_EMU_LONG_CHANNEL_DATA_C         : std_logic_vector(31 downto 0)    := x"00000000";           -- Long channel data for the TTC emulator
  constant REG_TTC_EMU_RESET_C                     : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register resets the TTC Emulator to the default state.
  constant REG_TTC_ECR_MONITOR_CLEAR_C             : std_logic_vector(64 downto 64)   := "0";                   -- Counts the number of ECRs received from the TTC system, any write to this register clears the counter
  constant REG_TTC_TTYPE_MONITOR_CLEAR_C           : std_logic_vector(64 downto 64)   := "0";                   -- Counts the number of TType received from the TTC system, any write to this register clears the counter
  constant REG_TTC_BCR_PERIODICITY_MONITOR_CLEAR_C : std_logic_vector(64 downto 64)   := "0";                   -- Counts the number of times the BCR period does not match 3564, any write to this register clears the counter
  constant REG_TTC_BCR_COUNTER_CLEAR_C             : std_logic_vector(64 downto 64)   := "0";                   -- Counts the number of times BCR is issued, any write to this register clears the counter
  constant REG_XOFF_FM_CH_FIFO_THRESH_LOW_C        : std_logic_vector(3 downto 0)     := x"b";                  -- Controls the low threshold of the channel fifo in FULL mode on which
                                                                                                                -- an Xon will be asserted, bitfields control 4 MSB
                                                                                                                
  constant REG_XOFF_FM_CH_FIFO_THRESH_HIGH_C       : std_logic_vector(3 downto 0)     := x"b";                  -- Controls the high threshold of the channel fifo in FULL mode on which
                                                                                                                -- an Xoff will be asserted, bitfields control 4 MSB
                                                                                                                
  constant REG_XOFF_FM_HIGH_THRESH_CLEAR_LATCH_C   : std_logic_vector(64 downto 64)   := "0";                   -- Writing this register will clear all CROSS_LATCHED bits
  constant REG_XOFF_FM_SOFT_XOFF_C                 : std_logic_vector(23 downto 0)    := x"000000";             -- Set any bit in this register to assert XOFF for the given channel, clearing bits will assert XON
  constant REG_XOFF_ENABLE_C                       : std_logic_vector(23 downto 0)    := x"000000";             -- Enable XOFF assertion (To Frontend) in case the FULL mode CH FIFO gets beyond thresholds. One bit per channel
  constant REG_DMA_BUSY_STATUS_CLEAR_LATCH_C       : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register clears TOHOST_BUSY_LATCHED
  constant REG_DMA_BUSY_STATUS_ENABLE_C            : std_logic_vector(4 downto 4)     := "0";                   -- Enable the DMA buffer on the server as a source of busy
  constant REG_FM_BUSY_CHANNEL_STATUS_CLEAR_LATCH_C: std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register will clear the BUSY_LATCHED bits
  constant REG_BUSY_MAIN_OUTPUT_FIFO_THRESH_BUSY_ENABLE_C: std_logic_vector(24 downto 24)   := "0";                   -- Enable busy generation if thresholds are crossed
  constant REG_BUSY_MAIN_OUTPUT_FIFO_THRESH_LOW_C  : std_logic_vector(23 downto 12)   := x"3ff";                -- Low, Negate threshold of busy generation from main output fifo
  constant REG_BUSY_MAIN_OUTPUT_FIFO_THRESH_HIGH_C : std_logic_vector(11 downto 0)    := x"4ff";                -- High, Assert threshold of busy generation from main output fifo
  constant REG_BUSY_MAIN_OUTPUT_FIFO_STATUS_CLEAR_LATCHED_C: std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register will clear the
  constant REG_ELINK_BUSY_ENABLE00_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE01_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE02_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE03_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE04_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE05_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE06_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE07_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE08_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE09_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE10_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE11_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE12_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE13_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE14_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE15_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE16_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE17_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE18_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE19_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE20_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE21_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE22_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_ELINK_BUSY_ENABLE23_C               : std_logic_vector(56 downto 0)    := "000000000000000000000000000000000000000000000000000000000"; -- Per elink (and FULL mode link) enable of the busy signal towards the LEMO output
  constant REG_BUSY_TOHOST_ENABLE_C                : std_logic_vector(0 downto 0)     := "0";                   -- Enable the busy ToHost Virtual Elink
  constant REG_HK_CTRL_I2C_CONFIG_TRIG_C           : std_logic_vector(1 downto 1)     := "0";                   -- i2c_config_trig
  constant REG_HK_CTRL_I2C_CLKFREQ_SEL_C           : std_logic_vector(0 downto 0)     := "0";                   -- i2c_clkfreq_sel
  constant REG_HK_CTRL_FMC_SI5345_INSEL_C          : std_logic_vector(6 downto 5)     := "00";                  -- Selects the input clock source
                                                                                                                --   0 : FPGA (FMC LA01)
                                                                                                                --   1 : FMC OSC (40.079 MHz)
                                                                                                                --   2 : FPGA (FMC LA18)
                                                                                                                
  constant REG_HK_CTRL_FMC_SI5345_A_C              : std_logic_vector(4 downto 3)     := "00";                  -- Si5345 I2C address select 2 LSB (0x0:default, dev id 0x68)
  constant REG_HK_CTRL_FMC_SI5345_OE_C             : std_logic_vector(2 downto 2)     := "1";                   -- Si5345 active low output enable  (0:enable)
  constant REG_HK_CTRL_FMC_SI5345_RSTN_C           : std_logic_vector(1 downto 1)     := "0";                   -- Si5345 active low output enable  (0:reset)
  constant REG_HK_CTRL_FMC_SI5345_SEL_C            : std_logic_vector(0 downto 0)     := "1";                   -- Si5345 programming mode
                                                                                                                --   1 : I2C mode (default)
                                                                                                                --   0 : SPI mode
                                                                                                                
  constant REG_HK_MON_FMC_SI5345_LOL_C             : std_logic_vector(1 downto 1)     := "0";                   -- Si5345 Loss Of Lock pin
  constant REG_HK_MON_FMC_SI5345_INTR_C            : std_logic_vector(0 downto 0)     := "0";                   -- Si5345 Interrupt flagging chip change of status
  constant REG_MMCM_MAIN_LCLK_SEL_C                : std_logic_vector(3 downto 3)     := "1";                   -- 1: LCLK
                                                                                                                -- 0: TTC
                                                                                                                
  constant REG_I2C_WR_I2C_WREN_C                   : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register triggers an I2C read or write sequence
  constant REG_I2C_WR_WRITE_2BYTES_C               : std_logic_vector(24 downto 24)   := "0";                   -- Write two bytes
  constant REG_I2C_WR_DATA_BYTE2_C                 : std_logic_vector(23 downto 16)   := x"00";                 -- Data byte 2
  constant REG_I2C_WR_DATA_BYTE1_C                 : std_logic_vector(15 downto 8)    := x"00";                 -- Data byte 1
  constant REG_I2C_WR_SLAVE_ADDRESS_C              : std_logic_vector(7 downto 1)     := "0000000";             -- Slave address
  constant REG_I2C_WR_READ_NOT_WRITE_C             : std_logic_vector(0 downto 0)     := "0";                   -- READ/<o>WRITE</o>
  constant REG_I2C_RD_I2C_RDEN_C                   : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register pops the last I2C data from the FIFO
  constant REG_INT_TEST_TRIGGER_C                  : std_logic_vector(64 downto 64)   := "0";                   -- Fire a test MSIx interrupt set in IRQ
  constant REG_INT_TEST_IRQ_C                      : std_logic_vector(3 downto 0)     := x"0";                  -- Set this field to a value equal to the MSIX interrupt to be fired. The write triggers the interrupt immediately.
  constant REG_CONFIG_FLASH_WR_FAST_WRITE_C        : std_logic_vector(57 downto 57)   := "0";                   -- Write command only. Only used for fast programming.
  constant REG_CONFIG_FLASH_WR_FAST_READ_C         : std_logic_vector(56 downto 56)   := "0";                   -- Status reading without command writing. Only used for fast programming.
  constant REG_CONFIG_FLASH_WR_PAR_CTRL_C          : std_logic_vector(55 downto 55)   := "0";                   -- Choose use FW or uC to select the Flash partition. 1 FW | 0 uC.
  constant REG_CONFIG_FLASH_WR_PAR_WR_C            : std_logic_vector(54 downto 53)   := "00";                  -- Choose Flash partition. Valid when PAR_CTRL is 1.
  constant REG_CONFIG_FLASH_WR_FLASH_SEL_C         : std_logic_vector(52 downto 52)   := "0";                   -- 1 takes control over flash, 0 gives JTAG control over flash
  constant REG_CONFIG_FLASH_WR_DO_INIT_C           : std_logic_vector(51 downto 51)   := "0";                   -- Untested feature, don't use it yet.
  constant REG_CONFIG_FLASH_WR_DO_READSTATUS_C     : std_logic_vector(50 downto 50)   := "0";                   -- Reads status from flash
  constant REG_CONFIG_FLASH_WR_DO_CLEARSTATUS_C    : std_logic_vector(49 downto 49)   := "0";                   -- Clears status reading from flash, back to normal flash operation
  constant REG_CONFIG_FLASH_WR_DO_ERASEBLOCK_C     : std_logic_vector(48 downto 48)   := "0";                   -- Erased the current block of the flash, this register has to be cleared by software
  constant REG_CONFIG_FLASH_WR_DO_UNLOCK_BLOCK_C   : std_logic_vector(47 downto 47)   := "0";                   -- Unlock writes to the current block, this register has to be cleared by software
  constant REG_CONFIG_FLASH_WR_DO_READ_C           : std_logic_vector(46 downto 46)   := "0";                   -- Reads the 16 bits from current address, this register has to be cleared by software
  constant REG_CONFIG_FLASH_WR_DO_WRITE_C          : std_logic_vector(45 downto 45)   := "0";                   -- Writes the 16 bits to current address, this register has to be cleared by software
  constant REG_CONFIG_FLASH_WR_DO_READDEVICEID_C   : std_logic_vector(44 downto 44)   := "0";                   -- DIN should return 0x0089, this register has to be cleared by software
  constant REG_CONFIG_FLASH_WR_DO_RESET_C          : std_logic_vector(43 downto 43)   := "0";                   -- Can be used in the future, currently disconnected in firmware
  constant REG_CONFIG_FLASH_WR_ADDRESS_C           : std_logic_vector(42 downto 16)   := "000000000000000000000000000"; -- Address for read and write operations (25 bits, upper 2 bits are controlled by uC)
  constant REG_CONFIG_FLASH_WR_WRITE_DATA_C        : std_logic_vector(15 downto 0)    := x"0000";               -- Value of data to write towards flash
  constant REG_RXUSRCLK_FREQ_CHANNEL_C             : std_logic_vector(37 downto 32)   := "000000";              -- Select the Transceiver channel to measure the clock from.
  constant REG_FELIG_L1ID_RESET_C                  : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register clears the FELIG L1ID
  constant REG_FELIG_DATA_GEN_CONFIG_00_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_00_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_00_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_00_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_00_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_00_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_01_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_01_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_01_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_01_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_01_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_01_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_02_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_02_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_02_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_02_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_02_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_02_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_03_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_03_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_03_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_03_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_03_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_03_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_04_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_04_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_04_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_04_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_04_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_04_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_05_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_05_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_05_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_05_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_05_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_05_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_06_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_06_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_06_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_06_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_06_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_06_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_07_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_07_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_07_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_07_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_07_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_07_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_08_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_08_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_08_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_08_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_08_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_08_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_09_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_09_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_09_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_09_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_09_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_09_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_10_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_10_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_10_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_10_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_10_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_10_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_11_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_11_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_11_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_11_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_11_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_11_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_12_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_12_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_12_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_12_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_12_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_12_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_13_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_13_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_13_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_13_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_13_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_13_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_14_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_14_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_14_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_14_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_14_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_14_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_15_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_15_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_15_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_15_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_15_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_15_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_16_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_16_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_16_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_16_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_16_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_16_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_17_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_17_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_17_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_17_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_17_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_17_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_18_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_18_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_18_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_18_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_18_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_18_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_19_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_19_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_19_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_19_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_19_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_19_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_20_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_20_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_20_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_20_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_20_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_20_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_21_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_21_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_21_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_21_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_21_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_21_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_22_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_22_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_22_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_22_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_22_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_22_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_DATA_GEN_CONFIG_23_USERDATA_C : std_logic_vector(63 downto 48)   := x"0000";               -- Sets static payload word. When PATTERN_SEL=1.
  constant REG_FELIG_DATA_GEN_CONFIG_23_CHUNK_LENGTH_C: std_logic_vector(47 downto 32)   := x"0000";               -- FELIG data generator chunk-length in bytes.
  constant REG_FELIG_DATA_GEN_CONFIG_23_RESET_C    : std_logic_vector(19 downto 15)   := "00000";               -- FELIG data generator reset. One bit per group, 0:normal operation, 1:egroup emulation held in reset.
  constant REG_FELIG_DATA_GEN_CONFIG_23_SW_BUSY_C  : std_logic_vector(14 downto 10)   := "00000";               -- FELIG elink bus state. One bit per group, 0:normal operation, 1:elink enter busy state.
  constant REG_FELIG_DATA_GEN_CONFIG_23_DATA_FORMAT_C: std_logic_vector(9 downto 5)     := "00000";               -- FELIG data generator format. 0:8b10b, 1:direct.
  constant REG_FELIG_DATA_GEN_CONFIG_23_PATTERN_SEL_C: std_logic_vector(4 downto 0)     := "00000";               -- FELIG data payload type. One bit per group, 0:byte counter, 1:USERDATA
  constant REG_FELIG_ELINK_CONFIG_00_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_00_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_00_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_01_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_01_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_01_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_02_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_02_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_02_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_03_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_03_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_03_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_04_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_04_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_04_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_05_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_05_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_05_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_06_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_06_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_06_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_07_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_07_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_07_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_08_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_08_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_08_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_09_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_09_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_09_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_10_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_10_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_10_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_11_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_11_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_11_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_12_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_12_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_12_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_13_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_13_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_13_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_14_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_14_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_14_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_15_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_15_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_15_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_16_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_16_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_16_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_17_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_17_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_17_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_18_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_18_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_18_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_19_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_19_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_19_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_20_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_20_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_20_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_21_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_21_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_21_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_22_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_22_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_22_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_CONFIG_23_ENDIAN_MOD_C  : std_logic_vector(39 downto 35)   := "00000";               -- FELIG elink data input endian control. One bit per egroup. 0:little-endian (8b10b), 1:big-endian.
  constant REG_FELIG_ELINK_CONFIG_23_INPUT_WIDTH_C : std_logic_vector(34 downto 30)   := "00000";               -- FELIG elink data input width. One bit per egroup. 0:8-bit (direct), 1:10-bit (8b10b).
  constant REG_FELIG_ELINK_CONFIG_23_OUTPUT_WIDTH_C: std_logic_vector(9 downto 0)     := "0000000000";          -- FELIG elink data output width.
  constant REG_FELIG_ELINK_ENABLE_00_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_01_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_02_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_03_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_04_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_05_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_06_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_07_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_08_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_09_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_10_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_11_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_12_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_13_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_14_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_15_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_16_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_17_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_18_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_19_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_20_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_21_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_22_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_ELINK_ENABLE_23_C             : std_logic_vector(39 downto 0)    := x"0000000000";         -- FELIG elink enable.  One bit per elink. 0:disabled, 1:enabled.
  constant REG_FELIG_GLOBAL_CONTROL_FAKE_L1A_RATE_C: std_logic_vector(63 downto 36)   := x"0000000";            -- Sets the internal fake L1 trigger rate. [25ns/LSB]
  constant REG_FELIG_GLOBAL_CONTROL_PICXO_OFFSET_PPM_C: std_logic_vector(35 downto 14)   := "0000000000000000000000"; -- When OFFSET_EN is 1, this directly sets the output frequency, within the given adjustment range.
  constant REG_FELIG_GLOBAL_CONTROL_TRACK_DATA_C   : std_logic_vector(12 downto 12)   := "0";                   -- FELIG GT core control.  Must be set to enable normal operation.
  constant REG_FELIG_GLOBAL_CONTROL_RXUSERRDY_C    : std_logic_vector(11 downto 11)   := "0";                   -- FELIG GT core control.  Must be set to enable normal operation.
  constant REG_FELIG_GLOBAL_CONTROL_TXUSERRDY_C    : std_logic_vector(10 downto 10)   := "0";                   -- FELIG GT core control.  Must be set to enable normal operation.
  constant REG_FELIG_GLOBAL_CONTROL_AUTO_RESET_C   : std_logic_vector(9 downto 9)     := "0";                   -- FELIG GT core control.  If set the GT core automatically resets on data error.
  constant REG_FELIG_GLOBAL_CONTROL_PICXO_RESET_C  : std_logic_vector(8 downto 8)     := "0";                   -- FELIG GT core control.  Manual PICXO reset.
  constant REG_FELIG_GLOBAL_CONTROL_GTTX_RESET_C   : std_logic_vector(7 downto 7)     := "0";                   -- FELIG GT core control.  Manual GT TX reset
  constant REG_FELIG_GLOBAL_CONTROL_CPLL_RESET_C   : std_logic_vector(6 downto 6)     := "0";                   -- FELIG GT core control.  Manual CPLL reset.
  constant REG_FELIG_GLOBAL_CONTROL_X3_X4_OUTPUT_SELECT_C: std_logic_vector(5 downto 0)     := "000000";              -- X3/X4 SMA output source select.
  constant REG_FELIG_LANE_CONFIG_00_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_00_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_00_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_00_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_00_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_00_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_00_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_00_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_00_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_00_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_00_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_01_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_01_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_01_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_01_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_01_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_01_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_01_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_01_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_01_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_01_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_01_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_02_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_02_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_02_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_02_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_02_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_02_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_02_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_02_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_02_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_02_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_02_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_03_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_03_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_03_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_03_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_03_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_03_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_03_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_03_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_03_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_03_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_03_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_04_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_04_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_04_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_04_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_04_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_04_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_04_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_04_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_04_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_04_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_04_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_05_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_05_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_05_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_05_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_05_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_05_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_05_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_05_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_05_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_05_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_05_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_06_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_06_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_06_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_06_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_06_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_06_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_06_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_06_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_06_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_06_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_06_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_07_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_07_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_07_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_07_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_07_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_07_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_07_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_07_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_07_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_07_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_07_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_08_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_08_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_08_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_08_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_08_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_08_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_08_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_08_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_08_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_08_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_08_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_09_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_09_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_09_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_09_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_09_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_09_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_09_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_09_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_09_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_09_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_09_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_10_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_10_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_10_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_10_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_10_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_10_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_10_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_10_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_10_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_10_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_10_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_11_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_11_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_11_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_11_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_11_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_11_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_11_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_11_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_11_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_11_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_11_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_12_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_12_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_12_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_12_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_12_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_12_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_12_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_12_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_12_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_12_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_12_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_13_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_13_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_13_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_13_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_13_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_13_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_13_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_13_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_13_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_13_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_13_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_14_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_14_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_14_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_14_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_14_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_14_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_14_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_14_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_14_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_14_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_14_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_15_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_15_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_15_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_15_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_15_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_15_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_15_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_15_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_15_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_15_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_15_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_16_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_16_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_16_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_16_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_16_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_16_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_16_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_16_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_16_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_16_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_16_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_17_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_17_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_17_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_17_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_17_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_17_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_17_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_17_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_17_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_17_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_17_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_18_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_18_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_18_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_18_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_18_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_18_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_18_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_18_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_18_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_18_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_18_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_19_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_19_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_19_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_19_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_19_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_19_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_19_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_19_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_19_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_19_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_19_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_20_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_20_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_20_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_20_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_20_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_20_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_20_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_20_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_20_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_20_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_20_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_21_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_21_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_21_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_21_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_21_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_21_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_21_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_21_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_21_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_21_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_21_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_22_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_22_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_22_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_22_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_22_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_22_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_22_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_22_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_22_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_22_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_22_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_LANE_CONFIG_23_B_CH_BIT_SEL_C : std_logic_vector(63 downto 42)   := "0000000000000000000000"; -- When OFFSET_EN is 1. this directly sets the output frequency. within the given adjustment range.
  constant REG_FELIG_LANE_CONFIG_23_A_CH_BIT_SEL_C : std_logic_vector(41 downto 35)   := "0000000";             -- Selects the bit from the received FELIX data from which to extract the L1A.
  constant REG_FELIG_LANE_CONFIG_23_LB_FIFO_DELAY_C: std_logic_vector(34 downto 30)   := "00000";               -- When the GTH or GTB loopback is enabled, this controls the loopback latency in clock cycles.
  constant REG_FELIG_LANE_CONFIG_23_ELINK_SYNC_C   : std_logic_vector(7 downto 7)     := "0";                   -- When set, synchronizes the elink word boundaries.  Must be set back to 0 to resume normal operation.
  constant REG_FELIG_LANE_CONFIG_23_PICXO_OFFEST_EN_C: std_logic_vector(6 downto 6)     := "0";                   -- FELIG TX frequency override. 0:frequency tracking enabled, 1:TX frequency set by PICXO_OFFSET_PPM.
  constant REG_FELIG_LANE_CONFIG_23_PI_HOLD_C      : std_logic_vector(5 downto 5)     := "0";                   -- FELIG phase-interpolator hold. 0:frequency tracking enabled, 1:freeze TX frequency.
  constant REG_FELIG_LANE_CONFIG_23_GBT_LB_ENABLE_C: std_logic_vector(4 downto 4)     := "0";                   -- FELIG GBT direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_23_GBH_LB_ENABLE_C: std_logic_vector(3 downto 3)     := "0";                   -- FELIG GTH direct loopback enable. 0:disabled, 1:enabled.
  constant REG_FELIG_LANE_CONFIG_23_L1A_SOURCE_C   : std_logic_vector(2 downto 2)     := "0";                   -- FELIG L1A data source select.  0:from local counter, 1:from FELIX.
  constant REG_FELIG_LANE_CONFIG_23_GBT_EMU_SOURCE_C: std_logic_vector(1 downto 1)     := "0";                   -- FELIG emulation data source select.  0:state-machine emulator, 1:ram-based emulator.
  constant REG_FELIG_LANE_CONFIG_23_FG_SOURCE_C    : std_logic_vector(0 downto 0)     := "0";                   -- FELIG link check data source selection control.  0:normal operation, 1:PRBS link checker (not elink emulation data)
  constant REG_FELIG_MON_FREQ_GLOBAL_XTAL_100MHZ_C : std_logic_vector(63 downto 32)   := x"00000000";           -- FELIG local oscillator frequency[Hz].
  constant REG_FELIG_MON_FREQ_GLOBAL_CLK_41_667MHZ_C: std_logic_vector(31 downto 0)    := x"00000000";           -- FELIG PCIE MGTREFCLK frequency[Hz].
  constant REG_FELIG_RESET_LB_FIFO_C               : std_logic_vector(63 downto 48)   := x"0000";               -- One bit per lane.  When set to 1, resets all loopback FIFOs.
  constant REG_FELIG_RESET_FRAMEGEN_C              : std_logic_vector(47 downto 24)   := x"000000";             -- One bit per lane.  When set to 1, resets all FELIG link checking logic.
  constant REG_FELIG_RESET_LANE_C                  : std_logic_vector(23 downto 0)    := x"000000";             -- One bit per lane.  When set to 1, resets all FELIG lane logic.
  constant REG_FELIG_RX_SLIDE_RESET_C              : std_logic_vector(23 downto 0)    := x"000000";             -- One bit per lane.  When set to 1, resets the gbt rx slide counter.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_00_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_00_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_01_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_01_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_02_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_02_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_03_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_03_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_04_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_04_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_05_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_05_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_06_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_06_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_07_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_07_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_08_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_08_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_09_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_09_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_10_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_10_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_11_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_11_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_12_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_12_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_13_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_13_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_14_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_14_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_15_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_15_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_16_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_16_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_17_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_17_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_18_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_18_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_19_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_19_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_20_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_20_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_21_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_21_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_22_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_22_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_23_ITKS_FIFO_CTL_C: std_logic_vector(19 downto 17)   := "000";                 -- data fifo control 2:rst 1:rd 0:wr.
  constant REG_FELIG_ITK_STRIPS_DATA_GEN_CONFIG_23_ITKS_FIFO_DATA_C: std_logic_vector(16 downto 0)    := "00000000000000000";   -- itks emu data 16:last word 15-0:data word
  constant REG_FMEMU_COUNTERS_WORD_CNT_C           : std_logic_vector(63 downto 48)   := x"0020";               -- Number of 32b words in one chunk
  constant REG_FMEMU_COUNTERS_IDLE_CNT_C           : std_logic_vector(47 downto 32)   := x"0003";               -- Minimum number of idles between chunks
  constant REG_FMEMU_COUNTERS_L1A_CNT_C            : std_logic_vector(31 downto 16)   := x"0100";               -- Number of chunks to send if not in TTC mode
  constant REG_FMEMU_COUNTERS_BUSY_TH_HIGH_C       : std_logic_vector(15 downto 8)    := x"14";                 -- Assert BUSY-ON above this threshold
  constant REG_FMEMU_COUNTERS_BUSY_TH_LOW_C        : std_logic_vector(7 downto 0)     := x"0f";                 -- De-assert BUSY-ON below this threshold
  constant REG_FMEMU_CONTROL_L1A_BITNR_C           : std_logic_vector(63 downto 56)   := x"30";                 -- Bitfield for L1A in TTC frame
  constant REG_FMEMU_CONTROL_XONXOFF_BITNR_C       : std_logic_vector(55 downto 48)   := x"20";                 -- Bitfield for Xon/Xoff in TTC frame
  constant REG_FMEMU_CONTROL_EMU_START_C           : std_logic_vector(47 downto 47)   := "0";                   -- Start emulator functionality
  constant REG_FMEMU_CONTROL_TTC_MODE_C            : std_logic_vector(46 downto 46)   := "0";                   -- Control the emulator by TTC input or by RegMap (1/0)
  constant REG_FMEMU_CONTROL_XONXOFF_C             : std_logic_vector(45 downto 45)   := "1";                   -- Enable Xon/Xoff functionality (1/0)
  constant REG_FMEMU_CONTROL_INLC_CRC32_C          : std_logic_vector(44 downto 44)   := "0";                   -- 0: No checksum
                                                                                                                -- 1: Append the data with a CRC32
                                                                                                                
  constant REG_FMEMU_CONTROL_BCR_C                 : std_logic_vector(43 downto 43)   := "0";                   -- Reset BCID to 0
  constant REG_FMEMU_CONTROL_ECR_C                 : std_logic_vector(42 downto 42)   := "0";                   -- Reset L1ID to 0
  constant REG_FMEMU_CONTROL_CONSTANT_CHUNK_LENGTH_C: std_logic_vector(41 downto 41)   := "0";                   -- Data source select
                                                                                                                -- 0: Random chunk length
                                                                                                                -- 1: Constant chunk length
                                                                                                                
  constant REG_FMEMU_CONTROL_FFU_FM_EMU_T_C        : std_logic_vector(16 downto 16)   := "0";                   -- For Future Use (trigger registers)
  constant REG_FMEMU_CONTROL_FE_BUSY_ENABLE_C      : std_logic_vector(0 downto 0)     := "1";                   -- Enable the BUSY mechanism if L1A counter passes threshold
  constant REG_FMEMU_RANDOM_RAM_ADDR_C             : std_logic_vector(9 downto 0)     := "0000000000";          -- Controls the address of the ramblock for the random number generator
  constant REG_FMEMU_RANDOM_RAM_WE_C               : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register (DATA) triggers a write to the ramblock
  constant REG_FMEMU_RANDOM_RAM_CHANNEL_SELECT_C   : std_logic_vector(39 downto 16)   := x"000000";             -- Enable write enable only for the selected channel
  constant REG_FMEMU_RANDOM_RAM_DATA_C             : std_logic_vector(15 downto 0)    := x"0000";               -- DATA field to be written to FMEMU_RANDOM_RAM_ADDR
  constant REG_FMEMU_RANDOM_CONTROL_SELECT_RANDOM_C: std_logic_vector(20 downto 20)   := "0";                   -- 1 enables the random chunk length, 0 uses a constant chunk length
  constant REG_FMEMU_RANDOM_CONTROL_SEED_C         : std_logic_vector(19 downto 10)   := "1000000000";          -- Seed for the random number generator, should not be 0
  constant REG_FMEMU_RANDOM_CONTROL_POLYNOMIAL_C   : std_logic_vector(9 downto 0)     := "1001000000";          -- POLYNOMIAL for the random number generator (10b LFSR) Bit9 should always be 1
  constant REG_FMEMU_CONFIG_WRADDR_C               : std_logic_vector(9 downto 0)     := "0000000000";          -- write enable for the FMEmu ram block
  constant REG_FMEMU_CONFIG_WE_C                   : std_logic_vector(64 downto 64)   := "0";                   -- Any write to register WRDATA triggers a write to the ramblock
  constant REG_FMEMU_CONFIG_CHANNEL_SELECT_C       : std_logic_vector(55 downto 32)   := x"000000";             -- Enable write enable only for the selected channel
  constant REG_FMEMU_CONFIG_WRDATA_C               : std_logic_vector(31 downto 0)    := x"00000000";           -- DATA field to be written to FMEMU_RANDOM_RAM_ADDR
  constant REG_WISHBONE_CONTROL_WRITE_NOT_READ_C   : std_logic_vector(32 downto 32)   := "0";                   -- wishbone write command wishbone read command
  constant REG_WISHBONE_CONTROL_ADDRESS_C          : std_logic_vector(31 downto 0)    := x"00000000";           -- Slave address for Wishbone bus
  constant REG_WISHBONE_WRITE_WRITE_ENABLE_C       : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register triggers a write to the Wupper to Wishbone fifo
  constant REG_WISHBONE_WRITE_DATA_C               : std_logic_vector(31 downto 0)    := x"00000000";           -- Wishbone
  constant REG_WISHBONE_READ_READ_ENABLE_C         : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register triggers a read from the Wishbone to Wupper fifo
  constant REG_IPBUS_WRITE_ADDRESS_C               : std_logic_vector(31 downto 0)    := x"00000000";           -- Address of the IPBus Write RAM
  constant REG_IPBUS_WRITE_DATA_WRITE_ENABLE_C     : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register triggers a write to the Wupper to IPBus inout RAM
  constant REG_IPBUS_WRITE_DATA_DATA_C             : std_logic_vector(63 downto 0)    := x"0000000000000000";   -- IPbus data to write to RAM
  constant REG_IPBUS_READ_ADDRESS_C                : std_logic_vector(31 downto 0)    := x"00000000";           -- Address of the IPBus Read RAM
  constant REG_GLOBAL_STRIPS_CONFIG_TEST_MODULE_MASK_C: std_logic_vector(63 downto 59)   := "00000";               -- (for tests only) contains R3 mask for the simulated trigger data
  constant REG_GLOBAL_STRIPS_CONFIG_TEST_R3L1_TAG_C: std_logic_vector(58 downto 52)   := "0000000";             -- (for tests only) contains R3 or L1 tag for the simulated trigger data
  constant REG_GLOBAL_STRIPS_CONFIG_TTC_GENERATE_GATING_ENABLE_C: std_logic_vector(51 downto 51)   := "0";                   -- Global control for gating signal generation. Enables generating trickle gating signal in response to TTC BCR. TRICKLE_TRIG_RUN must also be enabled for the trickle configuration to work. (See also BC_START, and BC_STOP fields)
  constant REG_GLOBAL_STRIPS_CONFIG_TTC_GATING_OVERRIDE_C: std_logic_vector(50 downto 50)   := "0";                   -- Overrides and disables gating signal generation when set to '1' (use if the elink is deadlocked and commands don't reach it).
  constant REG_GLOBAL_STRIPS_CONFIG_INVERT_AMAC_IN_C: std_logic_vector(4 downto 4)     := "0";                   -- Invert the polarity of all FELIX AMAC_IN elinks
  constant REG_GLOBAL_STRIPS_CONFIG_INVERT_AMAC_OUT_C: std_logic_vector(3 downto 3)     := "0";                   -- Invert the polarity of all FELIX AMAC_OUT elinks
  constant REG_GLOBAL_STRIPS_CONFIG_INVERT_DIN_C   : std_logic_vector(2 downto 2)     := "0";                   -- Invert the polarity of all FELIX 8-bit IN 8b10b elinks
  constant REG_GLOBAL_STRIPS_CONFIG_INVERT_R3L1_OUT_C: std_logic_vector(1 downto 1)     := "0";                   -- Invert the polarity of all FELIX R3L1 elinks
  constant REG_GLOBAL_STRIPS_CONFIG_INVERT_LCB_OUT_C: std_logic_vector(0 downto 0)     := "0";                   -- Invert the polarity of all FELIX LCB elinks
  constant REG_GLOBAL_TRICKLE_TRIGGER_C            : std_logic_vector(64 downto 64)   := "0";                   -- writing to this register issues a single trickle trigger for every LCB link connected to this FELIX device
  constant REG_STRIPS_R3_TRIGGER_C                 : std_logic_vector(64 downto 64)   := "0";                   -- (for tests only) simulate R3 trigger (issues 4-5 sequential triggers)
  constant REG_STRIPS_L1_TRIGGER_C                 : std_logic_vector(64 downto 64)   := "0";                   -- (for tests only) simulate L1 trigger (issues 4-5 sequential triggers)
  constant REG_STRIPS_R3L1_TRIGGER_C               : std_logic_vector(64 downto 64)   := "0";                   -- (for tests only) simulate simultaneous R3 and L1 trigger (issues 4-5 sequential triggers)
  constant REG_MROD_CTRL_OPTIONS_C                 : std_logic_vector(15 downto 8)    := x"00";                 -- Extra options for MROD
  constant REG_MROD_CTRL_ENASPARE1_C               : std_logic_vector(7 downto 7)     := "0";                   -- Enable spare1
  constant REG_MROD_CTRL_ENAMANSLIDE_C             : std_logic_vector(6 downto 6)     := "0";                   -- Enable Manual Slide in Rx Locking
  constant REG_MROD_CTRL_ENAPASSALL_C              : std_logic_vector(5 downto 5)     := "0";                   -- Enable PassAll in EmptySuppress
  constant REG_MROD_CTRL_ENATXCOUNT_C              : std_logic_vector(4 downto 4)     := "0";                   -- Enable SimpleCount in TxDriver for locking
  constant REG_MROD_CTRL_GOLTESTMODE_C             : std_logic_vector(3 downto 0)     := x"0";                  -- GOL Test Mode (emulate CSM):
                                                                                                                --   0: Run Data Emulator when 1;     0: stop, load emulator fifo
                                                                                                                --   1: Enable Circulate  when 1;     0: send fifo data only once
                                                                                                                --   2: Enable Triggered Mode when 1; 0: run continueously (no TTC)
                                                                                                                --   3: Enable pattern generator
                                                                                                                
  constant REG_MROD_TCVRCTRL_SLIDEMAX_C            : std_logic_vector(23 downto 16)   := x"ff";                 -- Maximum RXSLIDES before fire a TCVR reset
  constant REG_MROD_TCVRCTRL_SLIDEWAIT_C           : std_logic_vector(15 downto 8)    := x"20";                 -- RXclk delay in TCVR for next RX_SLIDE operation
  constant REG_MROD_TCVRCTRL_FRAMESIZE_C           : std_logic_vector(7 downto 0)     := x"14";                 -- Number of 32 data words in 1 frame
  constant REG_MROD_EP0_CSMENABLE_C                : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 CSM Data Enable channel 23-0
  constant REG_MROD_EP0_EMPTYSUPPR_C               : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 Set Empty Suppression channel 23-0
  constant REG_MROD_EP0_HPTDCMODE_C                : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 Set HPTDC Mode channel 23-0
  constant REG_MROD_EP0_CLRFIFOS_C                 : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 Clear FIFOs channel 23-0
  constant REG_MROD_EP0_EMULOADENA_C               : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 Emulator Load Enable channel 23-0
  constant REG_MROD_EP0_TRXLOOPBACK_C              : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 Transceiver Loopback Enable channel 23-0
  constant REG_MROD_EP0_TXCVRRESET_C               : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 Transceiver Reset all channel 23-0
  constant REG_MROD_EP0_RXRESET_C                  : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 Receiver Reset channel 23-0
  constant REG_MROD_EP0_TXRESET_C                  : std_logic_vector(23 downto 0)    := x"000000";             -- EP0 Transmitter Reset channel 23-0
  constant REG_MROD_EP1_CSMENABLE_C                : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 CSM Data Enable channel 23-0
  constant REG_MROD_EP1_EMPTYSUPPR_C               : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 Set Empty Suppression channel 23-0
  constant REG_MROD_EP1_HPTDCMODE_C                : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 Set HPTDC Mode channel 23-0
  constant REG_MROD_EP1_CLRFIFOS_C                 : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 Clear FIFOs channel 23-0
  constant REG_MROD_EP1_EMULOADENA_C               : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 Emulator Load Enable channel 23-0
  constant REG_MROD_EP1_TRXLOOPBACK_C              : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 Transceiver Loopback Enable channel 23-0
  constant REG_MROD_EP1_TXCVRRESET_C               : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 Transceiver Reset all channel 23-0
  constant REG_MROD_EP1_RXRESET_C                  : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 Receiver Reset channel 23-0
  constant REG_MROD_EP1_TXRESET_C                  : std_logic_vector(23 downto 0)    := x"000000";             -- EP1 Transmitter Reset channel 23-0
  -----------------------------------
  ---- GENERATED code END #3 ##  ----
  -----------------------------------

  --!
  --! --> MONITOR: Read Only User Application Registers (Read by PCIe)
  ------------------------------------
  ---- ## GENERATED code BEGIN #4 ----
  ------------------------------------

--
-- GenericBoardInformation
--
  type bitfield_generic_constants_r_type is record
    INTERRUPTS                     : std_logic_vector(15 downto 8);   -- Number of Interrupts
    DESCRIPTORS                    : std_logic_vector(7 downto 0);    -- Number of Descriptors
  end record;
  type bitfield_include_egroup_r_type is record
    TOHOST_32                      : std_logic_vector(9 downto 9);    -- ToHost EPATH32 is included in this EGROUP
    FROMHOST_02                    : std_logic_vector(8 downto 8);    -- FromHost EPATH02 is included in this EGROUP
    FROMHOST_04                    : std_logic_vector(7 downto 7);    -- FromHost EPATH04 is included in this EGROUP
    FROMHOST_08                    : std_logic_vector(6 downto 6);    -- FromHost EPATH8 is included in this EGROUP
    FROMHOST_HDLC                  : std_logic_vector(5 downto 5);    -- FromHost HDLC is included in this EGROUP
    TOHOST_02                      : std_logic_vector(4 downto 4);    -- ToHost EPATH02 is included in this EGROUP
    TOHOST_04                      : std_logic_vector(3 downto 3);    -- ToHost EPATH04 is included in this EGROUP
    TOHOST_08                      : std_logic_vector(2 downto 2);    -- ToHost EPATH08 is included in this EGROUP
    TOHOST_16                      : std_logic_vector(1 downto 1);    -- ToHost EPATH16 is included in this EGROUP
    TOHOST_HDLC                    : std_logic_vector(0 downto 0);    -- ToHost HDLC is included in this EGROUP
  end record;
  --Array of registers
  type bitfield_include_egroup_r_array_type is array (0 to 6) of bitfield_include_egroup_r_type;
  type bitfield_cr_generics_r_type is record
    XOFF_INCLUDED                  : std_logic_vector(2 downto 2);    -- Xoff bits (usually full mode) can be generated by the FromHost Central Router
    DIRECT_MODE_INCLUDED           : std_logic_vector(1 downto 1);    -- Indicates that the Direct mode functionality was built in the Central Router
    FROM_HOST_INCLUDED             : std_logic_vector(0 downto 0);    -- Indicates that the From Host path of the Central router was included in the design
  end record;
  type bitfield_axi_streams_tohost_r_type is record
    IC_INDEX                       : std_logic_vector(23 downto 16);  -- The AXIs ID (EPath-ID) of the ToHost IC E-Link
    EC_INDEX                       : std_logic_vector(15 downto 8);   -- The AXIs ID (EPath-ID) of the ToHost EC E-Link
    NUMBER_OF_STREAMS              : std_logic_vector(7 downto 0);    -- Total number of AXIs IDs (EPath-IDs) per physical link ToHost
  end record;
  type bitfield_axi_streams_fromhost_r_type is record
    IC_INDEX                       : std_logic_vector(23 downto 16);  -- The AXIs ID (EPath-ID) of the FromHost IC E-Link
    EC_INDEX                       : std_logic_vector(15 downto 8);   -- The AXIs ID (EPath-ID) of the FromHost EC E-Link
    NUMBER_OF_STREAMS              : std_logic_vector(7 downto 0);    -- Total number of AXIs IDs (EPath-IDs) per physical link FromHost
  end record;

  -- GenericBoardInformation
  type register_map_gen_board_info_type is record
    REG_MAP_VERSION                : std_logic_vector(15 downto 0);   -- Register Map Version, 5.0 formatted as 0x0500
    BOARD_ID_TIMESTAMP             : std_logic_vector(39 downto 0);   -- Board ID Date / Time in BCD format YYMMDDhhmm
    GIT_COMMIT_TIME                : std_logic_vector(39 downto 0);   -- Board ID GIT Commit time of current revision, Date / Time in BCD format YYMMDDhhmm
    GIT_TAG                        : std_logic_vector(63 downto 0);   -- String containing the current GIT TAG
    GIT_COMMIT_NUMBER              : std_logic_vector(31 downto 0);   -- Number of GIT commits after current GIT_TAG
    GIT_HASH                       : std_logic_vector(31 downto 0);   -- Short GIT hash (32 bit)
    GENERIC_CONSTANTS              : bitfield_generic_constants_r_type;
    NUM_OF_CHANNELS                : std_logic_vector(7 downto 0);    -- Number of GBT or FULL mode Channels
    CARD_TYPE                      : std_logic_vector(63 downto 0);   -- Card Type:
                                                                      --   - 709 (0x2c5): FLX709, VC709
                                                                      --   - 710 (0x2c6): FLX710, HTG710
                                                                      --   - 711 (0x2c7): FLX711, BNL711
                                                                      --   - 712 (0x2c8): FLX712, BNL712
                                                                      --   - 128 (0x080): FLX128, VCU128
                                                                      --   - 180 (0x0B4): FLX180, VMK180
                                                                      --   - 181 (0x0B5): FLX181, BNL181
                                                                      --   - 182 (0x0B6): FLX182, BNL182
                                                                      
    GENERATE_GBT                   : std_logic_vector(0 downto 0);    -- 1 when the GBT Wrapper is included in the design
    OPTO_TRX_NUM                   : std_logic_vector(7 downto 0);    -- Number of optical transceivers in the design
    GENERATE_TTC_EMU               : std_logic_vector(1 downto 1);    -- 1 when TTC emulator is generated
    INCLUDE_EGROUP                 : bitfield_include_egroup_r_array_type;
    WIDE_MODE                      : std_logic_vector(0 downto 0);    -- GBT is configured in Wide mode
    FIRMWARE_MODE                  : std_logic_vector(3 downto 0);    -- 0: GBT mode
                                                                      -- 1: FULL mode
                                                                      -- 2: LTDB mode (GBT mode with only IC and TTC links)
                                                                      -- 3: FEI4 mode
                                                                      -- 4: ITK Pixel
                                                                      -- 5: ITK Strip
                                                                      -- 6: FELIG
                                                                      -- 7: FULL mode emulator
                                                                      -- 8: FELIX_MROD mode
                                                                      -- 9: lpGBT mode
                                                                      -- 10: 25G Interlaken
                                                                      --             
                                                                      
    GTREFCLK_SOURCE                : std_logic_vector(1 downto 0);    -- 0: Transceiver reference Clock source from Si5345
                                                                      -- 1: Transceiver reference Clock source from Si5324
                                                                      -- 2: Transceiver reference Clock from internal BUFG (GREFCLK)
                                                                      
    CR_GENERICS                    : bitfield_cr_generics_r_type;  
    BLOCKSIZE                      : std_logic_vector(15 downto 0);   -- Number of bytes in a block
    PCIE_ENDPOINT                  : std_logic_vector(0 downto 0);    -- Indicator of the PCIe endpoint on BNL71x cards with two endpoints. 0 or 1
    CHUNK_TRAILER_32B              : std_logic_vector(0 downto 0);    -- Indicator that the chunk trailer is in the new 32-bit format
    NUMBER_OF_PCIE_ENDPOINTS       : std_logic_vector(1 downto 0);    -- Number of PCIe endpoints on the card. The BNL71x cards have 2 endpoints
    AXI_STREAMS_TOHOST             : bitfield_axi_streams_tohost_r_type;
    AXI_STREAMS_FROMHOST           : bitfield_axi_streams_fromhost_r_type;
    FROMHOST_LENGTH_IS_5BIT        : std_logic_vector(0 downto 0);    -- Set to 1 if the firmware is using the new FromHost data format as described in FLX-1355
    FULLMODE_HALFRATE              : std_logic_vector(0 downto 0);    -- If set to 1 the FULL mode firmware is running at 4.8Gb instead of the default 9.6Gb
    SUPPORT_HDLC_DELAY             : std_logic_vector(0 downto 0);    -- The HDLC encoders can offload a 1us delay as described in FLX-1826
end record;
--
-- CRToHostControlsAndMonitors
--
  type bitfield_crtohost_fifo_status_r_type is record
    FULL                           : std_logic_vector(47 downto 24);  -- Every bit represents the full flag of a channel FIFO
    FULL_LATCHED                   : std_logic_vector(23 downto 0);   -- like FULL but a latched state, clear by writing to this register
  end record;
  type bitfield_crtohost_dma_descriptor_2_r_type is record
    DESCR_READ                     : std_logic_vector(13 downto 11);  -- Read back the value of the descriptor assigned to AXIS_ID
  end record;

  -- CRToHostControlsAndMonitors
  type register_map_crtohost_monitor_type is record
    MAX_TIMEOUT                    : std_logic_vector(31 downto 0);   -- Maximum allowed timeout value
    CRTOHOST_FIFO_STATUS           : bitfield_crtohost_fifo_status_r_type;
    CRTOHOST_DMA_DESCRIPTOR_2      : bitfield_crtohost_dma_descriptor_2_r_type;
end record;
--
-- CRFromHostControlsAndMonitors
--
  -- Bitfields of CRFromHostControlsAndMonitors
  type bitfield_crfromhost_fifo_status_r_type is record
    FULL                           : std_logic_vector(47 downto 24);  -- Every bit represents the full flag of a channel FIFO
    FULL_LATCHED                   : std_logic_vector(23 downto 0);   -- like FULL but a latched state, clear by writing to this register
  end record;

  -- CRFromHostControlsAndMonitors
  type register_map_crfromhost_monitor_type is record
    CRFROMHOST_FIFO_STATUS         : bitfield_crfromhost_fifo_status_r_type;
end record;
--
-- DecodingControlsAndMonitors
--
  --Array of registers (std_logic_vector)
  type bitfield_decoding_link_aligned_r_array_type is  array (0 to 23) of  std_logic_vector(57 downto 0);   -- Every bit corresponds to an E-link on one (lp)GBT or FULL-mode frame. For FULL mode only bit 0 is used
  type bitfield_decoding_egroup_ctrl_r_type is record
    EPATH_ALMOST_FULL              : std_logic_vector(58 downto 51);  -- FIFO full indication
  end record;
  --Array of registers
  type bitfield_decoding_egroup_ctrl_r_array_type is array (0 to 6) of bitfield_decoding_egroup_ctrl_r_type;
  --Two dimensional array of registers
  type bitfield_decoding_egroup_ctrl_r_2d_array_type is array (0 to 11) of bitfield_decoding_egroup_ctrl_r_array_type;
  type bitfield_mini_egroup_tohost_r_type is record
    AUX_ALMOST_FULL                : std_logic_vector(12 downto 12);  -- Indicator that the AUX path FIFO is almost full
    IC_ALMOST_FULL                 : std_logic_vector(9 downto 9);    -- Indicator that the IC path FIFO is almost full
    EC_ALMOST_FULL                 : std_logic_vector(6 downto 6);    -- Indicator that the EC path FIFO is almost full
  end record;
  --Array of registers
  type bitfield_mini_egroup_tohost_r_array_type is array (0 to 23) of bitfield_mini_egroup_tohost_r_type;
  type bitfield_yarr_debug_allegroup_tohost_r_type is record
    CNT_RX_PACKET                  : std_logic_vector(31 downto 0);   -- Count packets of a given value
  end record;
  --Array of registers
  type bitfield_yarr_debug_allegroup_tohost_r_array_type is array (0 to 11) of bitfield_yarr_debug_allegroup_tohost_r_type;
  type bitfield_decoding_link_cb_r_type is record
    DESKEWED                       : std_logic_vector(61 downto 4);   -- Every bit corresponds to an E-link on one (lp)GBT frame. 
                                                                      -- Register indicates whether the E-link has been de-skewed in the channel. 
                                                                      -- E-link are grouped in a channel according to CBOPT
                                                                      
  end record;
  --Array of registers
  type bitfield_decoding_link_cb_r_array_type is array (0 to 11) of bitfield_decoding_link_cb_r_type;

  -- DecodingControlsAndMonitors
  type register_map_decoding_monitor_type is record
    DECODING_LINK_ALIGNED          : bitfield_decoding_link_aligned_r_array_type;
    DECODING_EGROUP_CTRL           : bitfield_decoding_egroup_ctrl_r_2d_array_type;
    MINI_EGROUP_TOHOST             : bitfield_mini_egroup_tohost_r_array_type;
    YARR_DEBUG_ALLEGROUP_TOHOST    : bitfield_yarr_debug_allegroup_tohost_r_array_type;
    DECODING_LINK_CB               : bitfield_decoding_link_cb_r_array_type;
end record;
--
-- EncodingControlsAndMonitors
--
  -- Bitfields of EncodingControlsAndMonitors
  type bitfield_encoding_egroup_ctrl_r_type is record
    EPATH_ALMOST_FULL              : std_logic_vector(58 downto 51);  -- Indiator that the EPATH FIFO is almost full
  end record;
  --Array of registers
  type bitfield_encoding_egroup_ctrl_r_array_type is array (0 to 4) of bitfield_encoding_egroup_ctrl_r_type;
  --Two dimensional array of registers
  type bitfield_encoding_egroup_ctrl_r_2d_array_type is array (0 to 11) of bitfield_encoding_egroup_ctrl_r_array_type;
  type bitfield_mini_egroup_fromhost_r_type is record
    AUX_ALMOST_FULL                : std_logic_vector(12 downto 12);  -- Indicator that the AUX Path FIFO is almost full
    IC_ALMOST_FULL                 : std_logic_vector(9 downto 9);    -- Indicator that the IC Path FIFO is almost full
    EC_ALMOST_FULL                 : std_logic_vector(6 downto 6);    -- Indicator that the EC Path FIFO is almost full
  end record;
  --Array of registers
  type bitfield_mini_egroup_fromhost_r_array_type is array (0 to 23) of bitfield_mini_egroup_fromhost_r_type;
  type bitfield_yarr_debug_allegroup_fromhost1_r_type is record
    CNT_TRIG_CMD                   : std_logic_vector(47 downto 16);  -- Number of issued triggers via cmd
    ERR_GENCALTRIG_DLY             : std_logic_vector(15 downto 8);   -- Number of mismatches between CNT_GENCALTRIG_DLY and REF_DLY_GENCALTRIG
  end record;
  --Array of registers
  type bitfield_yarr_debug_allegroup_fromhost1_r_array_type is array (0 to 11) of bitfield_yarr_debug_allegroup_fromhost1_r_type;
  type bitfield_yarr_debug_allegroup_fromhost2_r_type is record
    CNT_CMD                        : std_logic_vector(47 downto 16);  -- Number of issued commands
  end record;
  --Array of registers
  type bitfield_yarr_debug_allegroup_fromhost2_r_array_type is array (0 to 11) of bitfield_yarr_debug_allegroup_fromhost2_r_type;

  -- EncodingControlsAndMonitors
  type register_map_encoding_monitor_type is record
    ENCODING_EGROUP_CTRL           : bitfield_encoding_egroup_ctrl_r_2d_array_type;
    MINI_EGROUP_FROMHOST           : bitfield_mini_egroup_fromhost_r_array_type;
    YARR_DEBUG_ALLEGROUP_FROMHOST1 : bitfield_yarr_debug_allegroup_fromhost1_r_array_type;
    YARR_DEBUG_ALLEGROUP_FROMHOST2 : bitfield_yarr_debug_allegroup_fromhost2_r_array_type;
end record;
--
-- FrontendEmulatorControlsAndMonitors
--
  -- Bitfields of FrontendEmulatorControlsAndMonitors
  type bitfield_fe_emu_read_r_type is record
    DATA                           : std_logic_vector(32 downto 0);   -- Read back ramblock at FE_EMU_CONFIG.WRADDR
  end record;

  -- FrontendEmulatorControlsAndMonitors
  type register_map_gbtemu_monitor_type is record
    FE_EMU_READ                    : bitfield_fe_emu_read_r_type;  
end record;
--
-- LinkWrapperMonitors
--
  -- Bitfields of LinkWrapperMonitors
  type bitfield_gbt_version_r_type is record
    DATE                           : std_logic_vector(63 downto 48);  -- Date
    GBT_VERSION                    : std_logic_vector(47 downto 32);  -- GBT Version
    GTH_IP_VERSION                 : std_logic_vector(31 downto 16);  -- GTH IP Version
    RESERVED                       : std_logic_vector(15 downto 3);   -- Reserved
    GTHREFCLK_SEL                  : std_logic_vector(2 downto 2);    -- GTHREFCLK SEL
    RX_CLK_SEL                     : std_logic_vector(1 downto 1);    -- RX CLK SEL
    PLL_SEL                        : std_logic_vector(0 downto 0);    -- PLL SEL
  end record;
  type bitfield_gbt_pll_lock_r_type is record
    QPLL_LOCK                      : std_logic_vector(59 downto 48);  -- QPLL LOCK [11:0]
    CPLL_LOCK                      : std_logic_vector(47 downto 0);   -- CPLL LOCK [47:0]
  end record;

  -- LinkWrapperMonitors
  type register_map_link_monitor_type is record
    GBT_VERSION                    : bitfield_gbt_version_r_type;  
    GBT_TXRESET_DONE               : std_logic_vector(47 downto 0);   -- TX Reset done [47:0]
    GBT_RXRESET_DONE               : std_logic_vector(47 downto 0);   -- RX Reset done [47:0]
    GBT_TXFSMRESET_DONE            : std_logic_vector(47 downto 0);   -- TX FSM Reset done [47:0]
    GBT_RXFSMRESET_DONE            : std_logic_vector(47 downto 0);   -- RX FSM Reset done [47:0]
    GBT_CPLL_FBCLK_LOST            : std_logic_vector(47 downto 0);   -- CPLL FBCLK LOST [47:0]
    GBT_PLL_LOCK                   : bitfield_gbt_pll_lock_r_type; 
    GBT_RXCDR_LOCK                 : std_logic_vector(47 downto 0);   -- RX CDR LOCK [47:0]
    GBT_CLK_SAMPLED                : std_logic_vector(47 downto 0);   -- clk sampled [47:0]
    GBT_RX_IS_HEADER               : std_logic_vector(47 downto 0);   -- RX IS HEADER [47:0]
    GBT_RX_IS_DATA                 : std_logic_vector(47 downto 0);   -- RX IS DATA [47:0]
    GBT_RX_HEADER_FOUND            : std_logic_vector(47 downto 0);   -- RX HEADER FOUND [47:0]
    GBT_ALIGNMENT_DONE             : std_logic_vector(47 downto 0);   -- RX ALIGNMENT DONE [47:0]
    GBT_OUT_MUX_STATUS             : std_logic_vector(47 downto 0);   -- GBT output mux status [47:0]
    GBT_ERROR                      : std_logic_vector(47 downto 0);   -- Error flags [47:0]
    GBT_GBT_TOPBOT_C               : std_logic_vector(47 downto 0);   -- TopBot_c [47:0]
    GBT_FM_RX_DISP_ERROR1          : std_logic_vector(47 downto 0);   -- Rx disparity error [47:0]
    GBT_FM_RX_DISP_ERROR2          : std_logic_vector(47 downto 0);   -- Rx disparity error [96:48]
    GBT_FM_RX_NOTINTABLE1          : std_logic_vector(47 downto 0);   -- Rx not in table [47:0]
    GBT_FM_RX_NOTINTABLE2          : std_logic_vector(47 downto 0);   -- Rx not in table [96:48]
end record;
--
-- TTCBUSYControlsAndMonitors
--
  -- Bitfields of TTCBUSYControlsAndMonitors
  type bitfield_ttc_dec_ctrl_r_type is record
    BUSY_OUTPUT_STATUS             : std_logic_vector(14 downto 14);  -- Actual status of the BUSY LEMO output signal
  end record;
  type bitfield_ttc_dec_mon_r_type is record
    TH_FF_COUNT                    : std_logic_vector(15 downto 5);   -- ToHostData Fifo counts
    TH_FF_FULL                     : std_logic_vector(4 downto 4);    -- ToHostData Fifo status 1:full 0:not full
    TH_FF_EMPTY                    : std_logic_vector(3 downto 3);    -- ToHostData Fifo status 1:empty 0:not empty
    TTC_BIT_ERR                    : std_logic_vector(2 downto 0);    -- double bit, single bit and comm error in TTC data
  end record;
  --Array of registers (std_logic_vector)
  type bitfield_ttc_busy_accepted_r_array_type is  array (0 to 23) of  std_logic_vector(56 downto 0);   -- busy has been asserted by the given ELINK. Reset by writing to TTC_BUSY_CLEAR
  type bitfield_ttc_emu_r_type is record
    FULL                           : std_logic_vector(2 downto 2);    -- TTC Emulator memory full indication
  end record;
  type bitfield_ttc_ecr_monitor_r_type is record
    VALUE                          : std_logic_vector(31 downto 0);   -- Counts the number of ECRs received from the TTC system, any write to this register clears the counter
  end record;
  type bitfield_ttc_ttype_monitor_r_type is record
    VALUE                          : std_logic_vector(31 downto 0);   -- Counts the number of TType received from the TTC system, any write to this register clears the counter
  end record;
  type bitfield_ttc_bcr_periodicity_monitor_r_type is record
    VALUE                          : std_logic_vector(31 downto 0);   -- Counts the number of times the BCR period does not match 3564, any write to this register clears the counter
  end record;
  type bitfield_ttc_bcr_counter_r_type is record
    VALUE                          : std_logic_vector(31 downto 0);   -- Counts the number of times BCR is issued, any write to this register clears the counter
  end record;

  -- TTCBUSYControlsAndMonitors
  type register_map_ttc_monitor_type is record
    TTC_DEC_CTRL                   : bitfield_ttc_dec_ctrl_r_type; 
    TTC_DEC_MON                    : bitfield_ttc_dec_mon_r_type;  
    TTC_BUSY_ACCEPTED              : bitfield_ttc_busy_accepted_r_array_type;
    TTC_EMU                        : bitfield_ttc_emu_r_type;      
    TTC_L1ID_MONITOR               : std_logic_vector(31 downto 0);   -- Monitor L1ID and XL1ID.
    TTC_ECR_MONITOR                : bitfield_ttc_ecr_monitor_r_type;
    TTC_TTYPE_MONITOR              : bitfield_ttc_ttype_monitor_r_type;
    TTC_BCR_PERIODICITY_MONITOR    : bitfield_ttc_bcr_periodicity_monitor_r_type;
    TTC_BCR_COUNTER                : bitfield_ttc_bcr_counter_r_type;
end record;
--
-- XOFF_BUSYControlsAndMonitors
--
  type bitfield_xoff_fm_high_thresh_r_type is record
    CROSS_LATCHED                  : std_logic_vector(47 downto 24);  -- FIFO filled beyond the high threshold, 1 latch bit per channel
    CROSSED                        : std_logic_vector(23 downto 0);   -- FIFO filled beyond the high threshold, 1 bit per channel
  end record;
  type bitfield_dma_busy_status_r_type is record
    TOHOST_BUSY_LATCHED            : std_logic_vector(3 downto 3);    -- A tohost descriptor has passed BUSY_THRESHOLD_ASSERT in the past, busy flag was set
    TOHOST_BUSY                    : std_logic_vector(0 downto 0);    -- A tohost descriptor passed BUSY_THRESHOLD_ASSERT, busy flag set
  end record;
  type bitfield_fm_busy_channel_status_r_type is record
    BUSY_LATCHED                   : std_logic_vector(47 downto 24);  -- one Indicates that the given FULL mode channel has received BUSY-ON
    BUSY                           : std_logic_vector(23 downto 0);   -- one Indicates that the given FULL mode channel is currently in BUSY state
  end record;
  type bitfield_busy_main_output_fifo_status_r_type is record
    HIGH_THRESH_CROSSED_LATCHED    : std_logic_vector(2 downto 2);    -- Main output fifo has been full beyond HIGH THRESHOLD, write to clear
    HIGH_THRESH_CROSSED            : std_logic_vector(1 downto 1);    -- Main output fifo is full beyond HIGH THRESHOLD
    LOW_THRESH_CROSSED             : std_logic_vector(0 downto 0);    -- Main output fifo is full beyond LOW THRESHOLD
  end record;
  --Array of registers (std_logic_vector)
  type bitfield_xoff_peak_duration_r_array_type is  array (0 to 23) of  std_logic_vector(63 downto 0);   -- Maximum occurred duration of XOFF on the given channel in 25ns bins since reset
  --Array of registers (std_logic_vector)
  type bitfield_xoff_total_duration_r_array_type is  array (0 to 23) of  std_logic_vector(63 downto 0);   -- Total occurred duration of XOFF on the given channel in 25ns bins, divide by number of Xoffs to calculate the average since reset
  --Array of registers (std_logic_vector)
  type bitfield_xoff_count_r_array_type is  array (0 to 23) of  std_logic_vector(63 downto 0);   -- Total number of XOFF events per channel that occurred since a reset.

  -- XOFF_BUSYControlsAndMonitors
  type register_map_xoff_monitor_type is record
    XOFF_FM_LOW_THRESH_CROSSED     : std_logic_vector(23 downto 0);   -- FIFO filled beyond the low threshold, 1 bit per channel
    XOFF_FM_HIGH_THRESH            : bitfield_xoff_fm_high_thresh_r_type;
    DMA_BUSY_STATUS                : bitfield_dma_busy_status_r_type;
    FM_BUSY_CHANNEL_STATUS         : bitfield_fm_busy_channel_status_r_type;
    BUSY_MAIN_OUTPUT_FIFO_STATUS   : bitfield_busy_main_output_fifo_status_r_type;
    XOFF_PEAK_DURATION             : bitfield_xoff_peak_duration_r_array_type;
    XOFF_TOTAL_DURATION            : bitfield_xoff_total_duration_r_array_type;
    XOFF_COUNT                     : bitfield_xoff_count_r_array_type;
end record;
--
-- HouseKeepingControlsAndMonitors
--
  -- Bitfields of HouseKeepingControlsAndMonitors
  type bitfield_hk_ctrl_fmc_r_type is record
    SI5345_LOL                     : std_logic_vector(7 downto 7);    -- Loss of lock pin, only connected on FLX711
  end record;
  type bitfield_mmcm_main_r_type is record
    MAIN_INPUT                     : std_logic_vector(2 downto 1);    -- Main MMCM Oscillator Input
                                                                      -- 2: LCLK fixed
                                                                      -- 1: TTC fixed
                                                                      -- 0: selectable
                                                                      
    PLL_LOCK                       : std_logic_vector(0 downto 0);    -- Main MMCM PLL Lock Status
  end record;
  type bitfield_i2c_wr_r_type is record
    I2C_FULL                       : std_logic_vector(25 downto 25);  -- I2C FIFO full
  end record;
  type bitfield_i2c_rd_r_type is record
    I2C_EMPTY                      : std_logic_vector(8 downto 8);    -- I2C FIFO Empty
    I2C_DOUT                       : std_logic_vector(7 downto 0);    -- I2C READ Data
  end record;
  type bitfield_config_flash_rd_r_type is record
    PAR_RD                         : std_logic_vector(19 downto 18);  -- Show which Flash partition is selected.
    FLASH_REQ_DONE                 : std_logic_vector(17 downto 17);  -- Request done
    FLASH_BUSY                     : std_logic_vector(16 downto 16);  -- Flash operation busy
    READ_DATA                      : std_logic_vector(15 downto 0);   -- Value of data read from flash
  end record;
  type bitfield_si5324_status_r_type is record
    LOL                            : std_logic_vector(15 downto 8);   -- Loss of Lock Si5324
    LOS                            : std_logic_vector(8 downto 0);    -- Loss of Signal Si5324
  end record;
  type bitfield_rxusrclk_freq_r_type is record
    VALID                          : std_logic_vector(38 downto 38);  -- Indicates that the frequency measurement is valid
    VAL                            : std_logic_vector(31 downto 0);   -- Frequency in Hz of the selected channel
  end record;

  -- HouseKeepingControlsAndMonitors
  type register_map_hk_monitor_type is record
    HK_CTRL_FMC                    : bitfield_hk_ctrl_fmc_r_type;  
    MMCM_MAIN                      : bitfield_mmcm_main_r_type;    
    LMK_LOCKED                     : std_logic_vector(0 downto 0);    -- LMK Chip on BNL-711 locked
    FPGA_CORE_TEMP                 : std_logic_vector(11 downto 0);   -- XADC temperature monitor for the FPGA CORE
                                                                      -- for FLX709, FLX710
                                                                      -- temp (C)= ((FPGA_CORE_TEMP* 503.975)/4096)-273.15
                                                                      -- for FLX711
                                                                      -- temp (C)= ((FPGA_CORE_TEMP* 502.9098)/4096)-273.8195
                                                                      
    FPGA_CORE_VCCINT               : std_logic_vector(11 downto 0);   -- XADC voltage measurement VCCINT = (FPGA_CORE_VCCINT *3.0)/4096
    FPGA_CORE_VCCAUX               : std_logic_vector(11 downto 0);   -- XADC voltage measurement VCCAUX = (FPGA_CORE_VCCAUX *3.0)/4096
    FPGA_CORE_VCCBRAM              : std_logic_vector(11 downto 0);   -- XADC voltage measurement VCCBRAM = (FPGA_CORE_VCCBRAM *3.0)/4096
    FPGA_DNA                       : std_logic_vector(63 downto 0);   -- Unique identifier of the FPGA
    I2C_WR                         : bitfield_i2c_wr_r_type;       
    I2C_RD                         : bitfield_i2c_rd_r_type;       
    CONFIG_FLASH_RD                : bitfield_config_flash_rd_r_type;
    SI5324_STATUS                  : bitfield_si5324_status_r_type;
    TACH_CNT                       : std_logic_vector(19 downto 0);   -- Readout of the Fan tachometer speed of the BNL712 board
    RXUSRCLK_FREQ                  : bitfield_rxusrclk_freq_r_type;
end record;
--
-- Generators
--
  -- Bitfields of Generators
  type bitfield_felig_mon_ttc_0_r_type is record
    L1ID                           : std_logic_vector(63 downto 40);  -- Live TTC data monitor.
    XL1ID                          : std_logic_vector(39 downto 32);  -- Live TTC data monitor.
    BCID                           : std_logic_vector(31 downto 20);  -- Live TTC data monitor.
    RESERVED0                      : std_logic_vector(19 downto 16);  -- Live TTC data monitor.
    LEN                            : std_logic_vector(15 downto 8);   -- Live TTC data monitor.
    FMT                            : std_logic_vector(7 downto 0);    -- Live TTC data monitor.
  end record;
  --Array of registers
  type bitfield_felig_mon_ttc_0_r_array_type is array (0 to 23) of bitfield_felig_mon_ttc_0_r_type;
  type bitfield_felig_mon_ttc_1_r_type is record
    RESERVED1                      : std_logic_vector(63 downto 48);  -- Live TTC data monitor.
    TRIGGER_TYPE                   : std_logic_vector(47 downto 32);  -- Live TTC data monitor.
    ORBIT                          : std_logic_vector(31 downto 0);   -- Live TTC data monitor.
  end record;
  --Array of registers
  type bitfield_felig_mon_ttc_1_r_array_type is array (0 to 23) of bitfield_felig_mon_ttc_1_r_type;
  type bitfield_felig_mon_counters_r_type is record
    SLIDE_COUNT                    : std_logic_vector(63 downto 32);  -- Counts the number of rx slides commanded by the GBT logic.  Should be static once a link is established.
    FC_ERROR_COUNT                 : std_logic_vector(31 downto 0);   -- When FG_DATA_SELECT is 1, this counter reports the number of detected data errors.
  end record;
  --Array of registers
  type bitfield_felig_mon_counters_r_array_type is array (0 to 23) of bitfield_felig_mon_counters_r_type;
  type bitfield_felig_mon_freq_r_type is record
    TX                             : std_logic_vector(63 downto 32);  -- FELIG regenerated TX clock frequency[Hz].
    RX                             : std_logic_vector(31 downto 0);   -- FELIG recovered RX clock frequency[Hz].
  end record;
  --Array of registers
  type bitfield_felig_mon_freq_r_array_type is array (0 to 23) of bitfield_felig_mon_freq_r_type;
  --Array of registers (std_logic_vector)
  type bitfield_felig_mon_l1a_id_r_array_type is  array (0 to 23) of  std_logic_vector(31 downto 0);   -- FELIG's last L1 ID.
  type bitfield_felig_mon_picxo_r_type is record
    VLOT                           : std_logic_vector(53 downto 32);  -- Value indicates TX clock (recovered RX clock)  to RX reference clock frequency offset.
    ERROR                          : std_logic_vector(20 downto 0);   -- Value indicates RX to TX frequency tracking error.
  end record;
  --Array of registers
  type bitfield_felig_mon_picxo_r_array_type is array (0 to 23) of bitfield_felig_mon_picxo_r_type;
  --Array of registers (std_logic_vector)
  type bitfield_felig_mon_itk_strips_r_array_type is  array (0 to 23) of  std_logic_vector(2 downto 0);    -- data fifo status 2:write done 1:full 0:empty.
  type bitfield_fmemu_event_info_r_type is record
    L1ID                           : std_logic_vector(63 downto 32);  -- 32b field to show L1ID
    BCID                           : std_logic_vector(31 downto 0);   -- 32b field to show BCID
  end record;
  type bitfield_fmemu_control_r_type is record
    INT_STATUS_EMU                 : std_logic_vector(40 downto 32);  -- Read internal status emulator
  end record;

  -- Generators
  type register_map_generators_type is record
    FELIG_MON_TTC_0                : bitfield_felig_mon_ttc_0_r_array_type;
    FELIG_MON_TTC_1                : bitfield_felig_mon_ttc_1_r_array_type;
    FELIG_MON_COUNTERS             : bitfield_felig_mon_counters_r_array_type;
    FELIG_MON_FREQ                 : bitfield_felig_mon_freq_r_array_type;
    FELIG_MON_L1A_ID               : bitfield_felig_mon_l1a_id_r_array_type;
    FELIG_MON_PICXO                : bitfield_felig_mon_picxo_r_array_type;
    FELIG_MON_ITK_STRIPS           : bitfield_felig_mon_itk_strips_r_array_type;
    FMEMU_EVENT_INFO               : bitfield_fmemu_event_info_r_type;
    FMEMU_CONTROL                  : bitfield_fmemu_control_r_type;
end record;
--
-- Wishbone
--
  -- Bitfields of Wishbone
  type bitfield_wishbone_write_r_type is record
    FULL                           : std_logic_vector(32 downto 32);  -- Wishbone
  end record;
  type bitfield_wishbone_read_r_type is record
    EMPTY                          : std_logic_vector(32 downto 32);  -- Indicates that the Wishbone to Wupper fifo is empty
    DATA                           : std_logic_vector(31 downto 0);   -- Wishbone read data
  end record;
  type bitfield_wishbone_status_r_type is record
    INT                            : std_logic_vector(4 downto 4);    -- interrupt
    RETRY                          : std_logic_vector(3 downto 3);    -- Interface is not ready to accept data cycle should be retried
    STALL                          : std_logic_vector(2 downto 2);    -- When pipelined mode slave can't accept additional transactions in its queue
    ACKNOWLEDGE                    : std_logic_vector(1 downto 1);    -- Indicates the termination of a normal bus cycle
    ERROR                          : std_logic_vector(0 downto 0);    -- Address not mapped by the crossbar
  end record;

  -- Wishbone
  type wishbone_monitor_type is record
    WISHBONE_WRITE                 : bitfield_wishbone_write_r_type;
    WISHBONE_READ                  : bitfield_wishbone_read_r_type;
    WISHBONE_STATUS                : bitfield_wishbone_status_r_type;
end record;
--
-- MRODmonitors
--

  -- MRODmonitors
  type regmap_mrod_monitor_type is record
    MROD_EP0_CSMH_EMPTY            : std_logic_vector(23 downto 0);   -- EP0 CSM Handler FIFO Empty 23-0
    MROD_EP0_CSMH_FULL             : std_logic_vector(23 downto 0);   -- EP0 CSM Handler FIFO Full 23-0
    MROD_EP0_RXALIGNBSY            : std_logic_vector(23 downto 0);   -- EP0 Receiver Aligned monitor 23-0
    MROD_EP0_RXRECDATA             : std_logic_vector(23 downto 0);   -- EP0 Receiver Data monitor 23-0
    MROD_EP0_RXRECIDLES            : std_logic_vector(23 downto 0);   -- EP0 Receiver Idle monitor 23-0
    MROD_EP0_TXLOCKED              : std_logic_vector(23 downto 0);   -- EP0 Transmitter Locked monitor 23-0
    MROD_EP1_CSMH_EMPTY            : std_logic_vector(23 downto 0);   -- EP1 CSM Handler FIFO Empty 23-0
    MROD_EP1_CSMH_FULL             : std_logic_vector(23 downto 0);   -- EP1 CSM Handler FIFO Full 23-0
    MROD_EP1_RXALIGNBSY            : std_logic_vector(23 downto 0);   -- EP1 Receiver Aligned monitor 23-0
    MROD_EP1_RXRECDATA             : std_logic_vector(23 downto 0);   -- EP1 Receiver Data monitor 23-0
    MROD_EP1_RXRECIDLES            : std_logic_vector(23 downto 0);   -- EP1 Receiver Idle monitor 23-0
    MROD_EP1_TXLOCKED              : std_logic_vector(23 downto 0);   -- EP1 Transmitter Locked monitor 23-0
end record;
--
-- IPBus
--

  -- IPBus
  type ipbus_monitor_type is record
    IPBUS_READ_DATA                : std_logic_vector(63 downto 0);   -- IPbus data from Read RAM
    IPBUS_PKT_DONE                 : std_logic_vector(0 downto 0);    -- IPbus packet ready to read
end record;
  

  -- Monitor interface toward the dma_control block
  type register_map_monitor_type is record
    register_map_gen_board_info  : register_map_gen_board_info_type;
    register_map_crtohost_monitor  : register_map_crtohost_monitor_type;
    register_map_crfromhost_monitor  : register_map_crfromhost_monitor_type;
    register_map_decoding_monitor  : register_map_decoding_monitor_type;
    register_map_encoding_monitor  : register_map_encoding_monitor_type;
    register_map_gbtemu_monitor  : register_map_gbtemu_monitor_type;
    register_map_link_monitor  : register_map_link_monitor_type;
    register_map_ttc_monitor  : register_map_ttc_monitor_type;
    register_map_xoff_monitor  : register_map_xoff_monitor_type;
    register_map_hk_monitor  : register_map_hk_monitor_type;
    register_map_generators  : register_map_generators_type;
    wishbone_monitor  : wishbone_monitor_type;
    regmap_mrod_monitor  : regmap_mrod_monitor_type;
    ipbus_monitor  : ipbus_monitor_type;
  end record;
  
  -- Constants for unused monitor records

  constant register_map_gen_board_info_c : register_map_gen_board_info_type := (
    REG_MAP_VERSION                => (others => '0'),
    BOARD_ID_TIMESTAMP             => (others => '0'),
    GIT_COMMIT_TIME                => (others => '0'),
    GIT_TAG                        => (others => '0'),
    GIT_COMMIT_NUMBER              => (others => '0'),
    GIT_HASH                       => (others => '0'),
    GENERIC_CONSTANTS              => (others => (others => '0')),
    NUM_OF_CHANNELS                => (others => '0'),
    CARD_TYPE                      => (others => '0'),
    GENERATE_GBT                   => (others => '0'),
    OPTO_TRX_NUM                   => (others => '0'),
    GENERATE_TTC_EMU               => (others => '0'),
    INCLUDE_EGROUP                 => (others => (others => (others => '0'))),
    WIDE_MODE                      => (others => '0'),
    FIRMWARE_MODE                  => (others => '0'),
    GTREFCLK_SOURCE                => (others => '0'),
    CR_GENERICS                    => (others => (others => '0')),
    BLOCKSIZE                      => (others => '0'),
    PCIE_ENDPOINT                  => (others => '0'),
    CHUNK_TRAILER_32B              => (others => '0'),
    NUMBER_OF_PCIE_ENDPOINTS       => (others => '0'),
    AXI_STREAMS_TOHOST             => (others => (others => '0')),
    AXI_STREAMS_FROMHOST           => (others => (others => '0')),
    FROMHOST_LENGTH_IS_5BIT        => (others => '0'),
    FULLMODE_HALFRATE              => (others => '0'),
    SUPPORT_HDLC_DELAY             => (others => '0')
  );

  constant register_map_crtohost_monitor_c : register_map_crtohost_monitor_type := (
    MAX_TIMEOUT                    => (others => '0'),
    CRTOHOST_FIFO_STATUS           => (others => (others => '0')),
    CRTOHOST_DMA_DESCRIPTOR_2      => (others => (others => '0'))
  );

  constant register_map_crfromhost_monitor_c : register_map_crfromhost_monitor_type := (
    CRFROMHOST_FIFO_STATUS         => (others => (others => '0'))
  );

  constant register_map_decoding_monitor_c : register_map_decoding_monitor_type := (
    DECODING_LINK_ALIGNED          => (others => (others => '0')),
    DECODING_EGROUP_CTRL           => (others => (others => (others => (others => '0')))),
    MINI_EGROUP_TOHOST             => (others => (others => (others => '0'))),
    YARR_DEBUG_ALLEGROUP_TOHOST    => (others => (others => (others => '0'))),
    DECODING_LINK_CB               => (others => (others => (others => '0')))
  );

  constant register_map_encoding_monitor_c : register_map_encoding_monitor_type := (
    ENCODING_EGROUP_CTRL           => (others => (others => (others => (others => '0')))),
    MINI_EGROUP_FROMHOST           => (others => (others => (others => '0'))),
    YARR_DEBUG_ALLEGROUP_FROMHOST1 => (others => (others => (others => '0'))),
    YARR_DEBUG_ALLEGROUP_FROMHOST2 => (others => (others => (others => '0')))
  );

  constant register_map_gbtemu_monitor_c : register_map_gbtemu_monitor_type := (
    FE_EMU_READ                    => (others => (others => '0'))
  );

  constant register_map_link_monitor_c : register_map_link_monitor_type := (
    GBT_VERSION                    => (others => (others => '0')),
    GBT_TXRESET_DONE               => (others => '0'),
    GBT_RXRESET_DONE               => (others => '0'),
    GBT_TXFSMRESET_DONE            => (others => '0'),
    GBT_RXFSMRESET_DONE            => (others => '0'),
    GBT_CPLL_FBCLK_LOST            => (others => '0'),
    GBT_PLL_LOCK                   => (others => (others => '0')),
    GBT_RXCDR_LOCK                 => (others => '0'),
    GBT_CLK_SAMPLED                => (others => '0'),
    GBT_RX_IS_HEADER               => (others => '0'),
    GBT_RX_IS_DATA                 => (others => '0'),
    GBT_RX_HEADER_FOUND            => (others => '0'),
    GBT_ALIGNMENT_DONE             => (others => '0'),
    GBT_OUT_MUX_STATUS             => (others => '0'),
    GBT_ERROR                      => (others => '0'),
    GBT_GBT_TOPBOT_C               => (others => '0'),
    GBT_FM_RX_DISP_ERROR1          => (others => '0'),
    GBT_FM_RX_DISP_ERROR2          => (others => '0'),
    GBT_FM_RX_NOTINTABLE1          => (others => '0'),
    GBT_FM_RX_NOTINTABLE2          => (others => '0')
  );

  constant register_map_ttc_monitor_c : register_map_ttc_monitor_type := (
    TTC_DEC_CTRL                   => (others => (others => '0')),
    TTC_DEC_MON                    => (others => (others => '0')),
    TTC_BUSY_ACCEPTED              => (others => (others => '0')),
    TTC_EMU                        => (others => (others => '0')),
    TTC_L1ID_MONITOR               => (others => '0'),
    TTC_ECR_MONITOR                => (others => (others => '0')),
    TTC_TTYPE_MONITOR              => (others => (others => '0')),
    TTC_BCR_PERIODICITY_MONITOR    => (others => (others => '0')),
    TTC_BCR_COUNTER                => (others => (others => '0'))
  );

  constant register_map_xoff_monitor_c : register_map_xoff_monitor_type := (
    XOFF_FM_LOW_THRESH_CROSSED     => (others => '0'),
    XOFF_FM_HIGH_THRESH            => (others => (others => '0')),
    DMA_BUSY_STATUS                => (others => (others => '0')),
    FM_BUSY_CHANNEL_STATUS         => (others => (others => '0')),
    BUSY_MAIN_OUTPUT_FIFO_STATUS   => (others => (others => '0')),
    XOFF_PEAK_DURATION             => (others => (others => '0')),
    XOFF_TOTAL_DURATION            => (others => (others => '0')),
    XOFF_COUNT                     => (others => (others => '0'))
  );

  constant register_map_hk_monitor_c : register_map_hk_monitor_type := (
    HK_CTRL_FMC                    => (others => (others => '0')),
    MMCM_MAIN                      => (others => (others => '0')),
    LMK_LOCKED                     => (others => '0'),
    FPGA_CORE_TEMP                 => (others => '0'),
    FPGA_CORE_VCCINT               => (others => '0'),
    FPGA_CORE_VCCAUX               => (others => '0'),
    FPGA_CORE_VCCBRAM              => (others => '0'),
    FPGA_DNA                       => (others => '0'),
    I2C_WR                         => (others => (others => '0')),
    I2C_RD                         => (others => (others => '0')),
    CONFIG_FLASH_RD                => (others => (others => '0')),
    SI5324_STATUS                  => (others => (others => '0')),
    TACH_CNT                       => (others => '0'),
    RXUSRCLK_FREQ                  => (others => (others => '0'))
  );

  constant register_map_generators_c : register_map_generators_type := (
    FELIG_MON_TTC_0                => (others => (others => (others => '0'))),
    FELIG_MON_TTC_1                => (others => (others => (others => '0'))),
    FELIG_MON_COUNTERS             => (others => (others => (others => '0'))),
    FELIG_MON_FREQ                 => (others => (others => (others => '0'))),
    FELIG_MON_L1A_ID               => (others => (others => '0')),
    FELIG_MON_PICXO                => (others => (others => (others => '0'))),
    FELIG_MON_ITK_STRIPS           => (others => (others => '0')),
    FMEMU_EVENT_INFO               => (others => (others => '0')),
    FMEMU_CONTROL                  => (others => (others => '0'))
  );

  constant wishbone_monitor_c : wishbone_monitor_type := (
    WISHBONE_WRITE                 => (others => (others => '0')),
    WISHBONE_READ                  => (others => (others => '0')),
    WISHBONE_STATUS                => (others => (others => '0'))
  );

  constant regmap_mrod_monitor_c : regmap_mrod_monitor_type := (
    MROD_EP0_CSMH_EMPTY            => (others => '0'),
    MROD_EP0_CSMH_FULL             => (others => '0'),
    MROD_EP0_RXALIGNBSY            => (others => '0'),
    MROD_EP0_RXRECDATA             => (others => '0'),
    MROD_EP0_RXRECIDLES            => (others => '0'),
    MROD_EP0_TXLOCKED              => (others => '0'),
    MROD_EP1_CSMH_EMPTY            => (others => '0'),
    MROD_EP1_CSMH_FULL             => (others => '0'),
    MROD_EP1_RXALIGNBSY            => (others => '0'),
    MROD_EP1_RXRECDATA             => (others => '0'),
    MROD_EP1_RXRECIDLES            => (others => '0'),
    MROD_EP1_TXLOCKED              => (others => '0')
  );

  constant ipbus_monitor_c : ipbus_monitor_type := (
    IPBUS_READ_DATA                => (others => '0'),
    IPBUS_PKT_DONE                 => (others => '0')
  );
  -----------------------------------
  ---- GENERATED code END #4 ##  ----
  -----------------------------------

end package pcie_package ;

package body pcie_package is
    function to_sl( A: std_logic_vector) return std_logic is
    begin
        return A(A'low);
    end function to_sl;
    
    function or_reduce(slv : in std_logic_vector) return std_logic is
      variable res_v : std_logic := '0';  -- Null slv vector will also return '0'
    begin
      for i in slv'range loop
        res_v := res_v or slv(i);
      end loop;
      return res_v;
    end function;
    
end pcie_package;
