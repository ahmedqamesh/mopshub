//
// Verilog Module mopshub_lib.EPROC_IN2_DEC8b10b
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 19:58:01 04/02/21
//
// using Mentor Graphics HDL Designer(TM) 2018.1 (Build 12)
//

`resetall
`timescale 1ns/10ps
module EPROC_IN2_DEC8b10b (
    input   wire           bitCLK,
    input   wire           bitCLKx2,
    input   wire           rst,
    input   wire           swap_inputbits,
    input   wire           thCR_REVERSE_10B,
    input   wire    [1:0]  edataIN,
    output   wire    [9:0]  dataOUT,
    output   wire    dataOUTrdy



);


// ### Please start your Verilog code here ### 

endmodule
