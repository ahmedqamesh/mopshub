//
// Verilog Module mopshub_lib.tb_fifo_to_2K_18bit_wide
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 13:52:37 03/01/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module tb_fifo_to_2K_18bit_wide ;
  
  parameter DATA_WIDTH=18;
  
  wire [DATA_WIDTH-1:0] dout;
  wire almost_full,full,empty;
  wire prog_full;
  
  reg rd_en,wr_en,rd_clk,wr_clk;
  reg rst;
  
  //reg           enable;
  reg tx_fifo_pfull;
  wire done;               // dbg
  wire [DATA_WIDTH-1:0] din_gen;
  wire wen; //wr_en signal

  
  
  fh_epath_fifo2K_18bit_wide fifo2K_18bit_wide(.dout(dout),
  .full(full),
  .empty(empty),
  .prog_full(prog_full),
  .almost_full(almost_full),
  .din(din_gen),
  .rd_en(rd_en),
  .wr_en(wen),
  .rd_clk(rd_clk),
  .wr_clk(wr_clk),
  .rst(rst));
  
  data_generator DataGEN(
  .clk_usr(wr_clk),
  .enable(~rst),
  .loop_en(~rst),
  .done(done),
  .tx_fifo_pfull(tx_fifo_pfull),
  .dout(din_gen),
  .wen(wen)
  ); 
  
  
  //initial #100 $stop;
  initial begin 
    rd_clk=0; 
    forever #1 rd_clk=~rd_clk; 
  end
  
  initial begin 
    wr_clk=0; 
    forever #1 wr_clk=~wr_clk; 
  end  
  
  
  initial 
  begin 
    rd_en= 0;
    wr_en= 0;
    tx_fifo_pfull = 0;
    rst=1;
    #2 rst=0;
    rd_en=1;
  end                     
endmodule