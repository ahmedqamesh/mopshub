//
// Verilog Module mopshub_lib.sys_clk_emci
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 19:02:03 03/18/22
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
//----------------------------------------------------------------------------
// User entered comments
//----------------------------------------------------------------------------
// None
//
//----------------------------------------------------------------------------
//  Output     Output      Phase    Duty Cycle   Pk-to-Pk     Phase
//   Clock     Freq (MHz)  (degrees)    (%)     Jitter (ps)  Error (ps)
//----------------------------------------------------------------------------
// __clk_40__40.00000______0.000______50.0______153.625_____95.014
// __clk_80__80.00000______0.000______50.0______132.221_____95.014
// __clk_tx__160.00000______0.000______50.0______116.326_____95.014
// __clk_rx__40.00000______0.000______50.0______153.625_____95.014
//
//----------------------------------------------------------------------------
// Input Clock   Freq (MHz)    Input Jitter (UI)
//----------------------------------------------------------------------------
// __primary__________80.000____________0.010
`resetall
`timescale 1ns/10ps
module ip_sys_clk_emci( 
  output        clk_40,
  output        clk_80,
  output        clk_tx,
  output        clk_rx,
  // Status and control signals
  output        locked,
  input         clk_in1_p,
  input         clk_in1_n
 );

  // Input buffering
  //------------------------------------
//wire clk_local_sig;
wire clk_in1_mopshub_emci_clk_wiz_0_0;
  IBUFDS clkin1_ibufds ////The IBUFGDS are used to connect an input buffer that can be connected to a BUFG.
   (.O  (clk_in1_mopshub_emci_clk_wiz_0_0),//(clk_local_sig),
    .I  (clk_in1_p),
    .IB (clk_in1_n));
    
//  BUFG clkin_buf 
//   (.O   (clk_in1_mopshub_emci_clk_wiz_0_0),
//    .I   (clk_local_sig));
//
//


  // Clocking PRIMITIVE
  //------------------------------------

  // Instantiation of the MMCM PRIMITIVE
  //    * Unused inputs are tied off
  //    * Unused outputs are labeled unused

  wire        clk_40_mopshub_emci_clk_wiz_0_0;
  wire        clk_80_mopshub_emci_clk_wiz_0_0;
  wire        clk_tx_mopshub_emci_clk_wiz_0_0;
  wire        clk_rx_mopshub_emci_clk_wiz_0_0;
  wire        clk_out5_mopshub_emci_clk_wiz_0_0;
  wire        clk_out6_mopshub_emci_clk_wiz_0_0;
  wire        clk_out7_mopshub_emci_clk_wiz_0_0;

  wire [15:0] do_unused;
  wire        drdy_unused;
  wire        psdone_unused;
  wire        locked_int;
  wire        clkfbout_mopshub_emci_clk_wiz_0_0;
  wire        clkfbout_buf_mopshub_emci_clk_wiz_0_0;
  wire        clkfboutb_unused;
    wire clkout0b_unused;
   wire clkout1b_unused;
   wire clkout2b_unused;
   wire clkout3b_unused;
   wire clkout4_unused;
  wire        clkout5_unused;
  wire        clkout6_unused;
  wire        clkfbstopped_unused;
  wire        clkinstopped_unused;


  
    MMCME4_ADV

  #(.BANDWIDTH            ("OPTIMIZED"),
    .CLKOUT4_CASCADE      ("FALSE"),
    .COMPENSATION         ("AUTO"),
    .STARTUP_WAIT         ("FALSE"),
    .DIVCLK_DIVIDE        (1),
    .CLKFBOUT_MULT_F      (14.000),
    .CLKFBOUT_PHASE       (0.000),
    .CLKFBOUT_USE_FINE_PS ("FALSE"),
    .CLKOUT0_DIVIDE_F     (28.000),
    .CLKOUT0_PHASE        (0.000),
    .CLKOUT0_DUTY_CYCLE   (0.500),
    .CLKOUT0_USE_FINE_PS  ("FALSE"),
    .CLKOUT1_DIVIDE       (14),
    .CLKOUT1_PHASE        (0.000),
    .CLKOUT1_DUTY_CYCLE   (0.500),
    .CLKOUT1_USE_FINE_PS  ("FALSE"),
    .CLKOUT2_DIVIDE       (7),
    .CLKOUT2_PHASE        (0.000),
    .CLKOUT2_DUTY_CYCLE   (0.500),
    .CLKOUT2_USE_FINE_PS  ("FALSE"),
    .CLKOUT3_DIVIDE       (28),
    .CLKOUT3_PHASE        (0.000),
    .CLKOUT3_DUTY_CYCLE   (0.500),
    .CLKOUT3_USE_FINE_PS  ("FALSE"),
    .CLKIN1_PERIOD        (12.500))
  
  mmcme4_adv_inst
    // Output clocks
   (
    .CLKFBOUT            (clkfbout_mopshub_emci_clk_wiz_0_0),
    .CLKFBOUTB           (clkfboutb_unused),
    .CLKOUT0             (clk_40_mopshub_emci_clk_wiz_0_0),
    .CLKOUT0B            (clkout0b_unused),
    .CLKOUT1             (clk_80_mopshub_emci_clk_wiz_0_0),
    .CLKOUT1B            (clkout1b_unused),
    .CLKOUT2             (clk_tx_mopshub_emci_clk_wiz_0_0),
    .CLKOUT2B            (clkout2b_unused),
    .CLKOUT3             (clk_rx_mopshub_emci_clk_wiz_0_0),
    .CLKOUT3B            (clkout3b_unused),
    .CLKOUT4             (clkout4_unused),
    .CLKOUT5             (clkout5_unused),
    .CLKOUT6             (clkout6_unused),
     // Input clock control
    .CLKFBIN             (clkfbout_buf_mopshub_emci_clk_wiz_0_0),
    .CLKIN1              (clk_in1_mopshub_emci_clk_wiz_0_0),
    .CLKIN2              (1'b0),
     // Tied to always select the primary input clock
    .CLKINSEL            (1'b1),
    // Ports for dynamic reconfiguration
    .DADDR               (7'h0),
    .DCLK                (1'b0),
    .DEN                 (1'b0),
    .DI                  (16'h0),
    .DO                  (do_unused),
    .DRDY                (drdy_unused),
    .DWE                 (1'b0),
    .CDDCDONE            (),
    .CDDCREQ             (1'b0),
    // Ports for dynamic phase shift
    .PSCLK               (1'b0),
    .PSEN                (1'b0),
    .PSINCDEC            (1'b0),
    .PSDONE              (psdone_unused),
    // Other control and status signals
    .LOCKED              (locked_int),
    .CLKINSTOPPED        (clkinstopped_unused),
    .CLKFBSTOPPED        (clkfbstopped_unused),
    .PWRDWN              (1'b0),
    .RST                 (1'b0));

  assign locked = locked_int;
// Clock Monitor clock assigning
//--------------------------------------
 // Output buffering
  //-----------------------------------

  BUFG clkf_buf
   (.O (clkfbout_buf_mopshub_emci_clk_wiz_0_0),
    .I (clkfbout_mopshub_emci_clk_wiz_0_0));

  BUFG clkout1_buf
   (.O   (clk_40),
    .I   (clk_40_mopshub_emci_clk_wiz_0_0));


  BUFG clkout2_buf
   (.O   (clk_80),
    .I   (clk_80_mopshub_emci_clk_wiz_0_0));

  BUFG clkout3_buf
   (.O   (clk_tx),
    .I   (clk_tx_mopshub_emci_clk_wiz_0_0));

  BUFG clkout4_buf
   (.O   (clk_rx),
    .I   (clk_rx_mopshub_emci_clk_wiz_0_0));



endmodule