//
// Verilog Module mopshub_lib.tb_FIFO_to_Elink
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 12:41:49 03/19/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module tb_FIFO_to_Elink ;
  parameter DATA_WIDTH=8;
  parameter DATA_OUT_WIDTH = 10;
  reg                            clk_160;
  reg                            rst; 
  wire                            clk_80;
  wire                            clk_40; 
  wire                            gen_clk;
  
  //FIFO_to_Elink Signals
  wire                         DATA1bitOUT; 
  wire    [1:0]                elink2bit; 
  
  //FIFO Signals
  wire [DATA_OUT_WIDTH-1:0] Dout;
  wire doutRdy;
  wire getDataTrig;
  //data Genrator Signal
  wire [DATA_WIDTH-1:0] GEN_EDATA_8bit;
  wire tx_fifo_pfull;
  wire wr_en; 
  wire [1:0]delimeter;
  wire done; 
  reg enable;
  
  //GBTX Emulator Signals
  wire [DATA_WIDTH-1:0] DEC_EDATA_OUT_8bit;
  wire [DATA_OUT_WIDTH-1:0] ENC_EDATA_OUT_10bit;
  wire ko;
  wire code_err;
  wire disp_err;
  
  assign Dout = MUT.efifoDout;
  assign doutRdy = MUT.doutRdy;
  assign getDataTrig = MUT.efifoRE;
  
  data_generator DataGEN(
  .clk_usr          (gen_clk),
  .enable           (enable),
  .loop_en          (enable),
  .done             (done),
  .tx_fifo_pfull    (tx_fifo_pfull),
  .dout             (GEN_EDATA_8bit),
  .delimeter        (delimeter),
  .wr_en            (wr_en)
  );
  
  FIFO_to_Elink MUT(
  .wr_clk          (clk_40),
  .clk_80           (clk_80),
  .bitCLKx4         (clk_160),
  .rst              (rst),
  .fifo_flush       (rst),
  .efifoWe          (wr_en),
  .efifoDin         ({delimeter,GEN_EDATA_8bit}),
  .efifoPfull       (tx_fifo_pfull),
  .DATA1bitOUT      (DATA1bitOUT),
  .elink2bit        (elink2bit)
  );
  
  
  GBTX_Emulator U_1( 
  .ko               (ko), 
  .code_err         (code_err), 
  .disp_err         (disp_err), 
  .rst              (rst), 
  .bitCLK           (clk_40),
  .dataout          (DEC_EDATA_OUT_8bit), 
  .enc10bit_out_sig (ENC_EDATA_OUT_10bit),
  .EDATA_2bit       (elink2bit),
  .datain_valid     (~rst),
  .data_10b_in      (), 
  .data_10b_en      ()
  );
  
  //clk_40 to FIFO //40 Mb 
  //Freq. clk_40 = Freq. clk_160 / 4 [=40 MHz]
  clock_divider #(4) div_0(
  .clock_in(clk_160),
  .clock_out(clk_40)//Equivalent to the bitCLK
  );
  
  //Generator clk
  //Freq. gen_clk = Freq. clk_160 / 4 [=40 MHz]
  clock_divider #(4) div_1(
  .clock_in(clk_160),
  .clock_out(gen_clk)//Equivalent to the clk_40
  );
  //Generator clk_80 // 80 Mb
  //Freq. clk_80 = Freq. clk_160 / 2 [=80 MHz]
  clock_divider #(2) div_2(
  .clock_in(clk_160),
  .clock_out(clk_80)//Equivalent to the bitCLKx2
  );
  
  initial begin 
    clk_160=0; 
    forever #1 clk_160=~clk_160; //Equivalent to the bitCLKx4
  end
  
  initial 
  begin 
    enable = 1;
    rst = 1;
    #1 rst =0;
  end 
  always@(done)
    begin
      enable =0;
      #16;
      enable =1;
    end
  
endmodule
