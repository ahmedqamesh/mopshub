//
// Verilog Module mopshub_lib.tb_FIFO_to_Elink
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 12:41:49 03/19/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module tb_FIFO_to_Elink ;
  parameter DATA_WIDTH=18;
  parameter DATA_OUT_WIDTH = 10;
  wire                            clk_80;
  wire                            wr_clk; 
  reg                            clk_160;
  wire                            gen_clk;
  reg                            rst; 
  //FIFO_to_Elink Signals
  wire                         DATA1bitOUT; 
  wire    [1:0]                elink2bit; 
  
  //FIFO Signals
  wire [DATA_OUT_WIDTH-1:0] Dout;
  wire doutRdy;
  wire getDataTrig;
  //data Genrator Signal
  
  wire done;          
  wire [DATA_WIDTH-1:0] GEN_EDATA_18bit;
  wire wen; //wr_en signal
  
  //GBTX Emulator Signals
  wire [7:0] DEC_EDATA_OUT_8bit;
  wire [9:0] ENC_EDATA_OUT_10bit;
  wire ko;
  wire code_err;
  wire disp_err;
  
  
  assign Dout = MUT.efifoDout;
  assign doutRdy = MUT.doutRdy;
  assign getDataTrig = MUT.efifoRE;
  
  data_generator DataGEN(
  .clk_usr          (gen_clk),
  .enable           (~rst),
  .loop_en          (~rst),
  .done             (done),
  .tx_fifo_pfull    (1'b0),
  .dout             (GEN_EDATA_18bit),
  .wen              (wen)
  );
  
  
  FIFO_to_Elink MUT(
  .wr_clk          (wr_clk),
  .clk_80           (clk_80),
  .bitCLKx4         (clk_160),
  .rst              (rst),
  .fifo_flush       (rst),
  .efifoWe          (wen),
  .efifoDin         (GEN_EDATA_18bit),
  .efifoPfull       (),
  .DATA1bitOUT      (DATA1bitOUT),
  .elink2bit        (elink2bit)
  );
  
  
  GBTX_Emulator U_1( 
  .ko               (ko), 
  .code_err         (code_err), 
  .disp_err         (disp_err), 
  .rst              (rst), 
  .bitCLK           (clk_80),
  .dataout          (DEC_EDATA_OUT_8bit), 
  .enc10bit_out_sig (ENC_EDATA_OUT_10bit),
  .EDATA_2bit       (elink2bit),
  .datain_valid     (~rst),
  .data_10b_in      (), 
  .data_10b_en      ()
  );
  
  //initial #5000 $stop;
  //Wr_clk to FIFO //40 Mb 
  //Freq. Wr_clk = Freq. rd_clk / 4 [=40 MHz]
  clock_divider #(4) div_0(
  .clock_in(clk_160),
  .clock_out(wr_clk)//Equivalent to the bitCLK
  );
  

  //Generator clk
  //Freq. gen_clk = Freq. rd_clk / 4 [=40 MHz]
  clock_divider #(4) div_1(
  .clock_in(clk_160),
  .clock_out(gen_clk)//Equivalent to the wr_clk
  );
  
  
  //Generator clk // 80 Mb
  //Freq. gen_clk = Freq. rd_clk / 4 [=40 MHz]
  clock_divider #(2) div_2(
  .clock_in(clk_160),
  .clock_out(clk_80)//Equivalent to the wr_clk
  );
  
  initial begin 
    clk_160=0; 
    forever #1 clk_160=~clk_160; 
  end

  initial 
  begin 
    //rst module
    rst = 1;
    #10 rst =0;
  end 
  
  
endmodule
