--! This file is part of the FELIX firmware distribution (https://gitlab.cern.ch/atlas-tdaq-felix/firmware/).
--! Copyright (C) 2001-2021 CERN for the benefit of the ATLAS collaboration.
--! Authors:
--!               Marius Wensing
--!               Nico Giangiacomi
--!               Frans Schreuder
--! 
--!   Licensed under the Apache License, Version 2.0 (the "License");
--!   you may not use this file except in compliance with the License.
--!   You may obtain a copy of the License at
--!
--!       http://www.apache.org/licenses/LICENSE-2.0
--!
--!   Unless required by applicable law or agreed to in writing, software
--!   distributed under the License is distributed on an "AS IS" BASIS,
--!   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--!   See the License for the specific language governing permissions and
--!   limitations under the License.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

--library XPM;
--use XPM.VCOMPONENTS.ALL;

use work.axi_stream_package.ALL;

entity Axis8Fifo is
	generic (
		DEPTH : integer;
		CLOCKING_MODE : string := "independent_clock";
		RELATED_CLOCKS : integer range 0 to 1 := 0;
		FIFO_MEMORY_TYPE : string := "auto";
		PACKET_FIFO : string := "false";
		USE_BUILT_IN_FIFO : std_logic := '1'
	);
	port (
		-- axi stream slave
		s_axis_aresetn : in std_logic;
		s_axis_aclk : in std_logic;
		s_axis : in axis_8_type;
		s_axis_tready : out std_logic;

		-- axi stream master
		m_axis_aclk : in std_logic;
		m_axis : out axis_8_type;
		m_axis_tready : in std_logic;
		almost_full : out std_logic
	);
end Axis8Fifo;

architecture rtl of Axis8Fifo is


COMPONENT axi8_fifo_bif
  PORT (
    wr_rst_busy : OUT STD_LOGIC;
    rd_rst_busy : OUT STD_LOGIC;
    m_aclk : IN STD_LOGIC;
    s_aclk : IN STD_LOGIC;
    s_aresetn : IN STD_LOGIC;
    s_axis_tvalid : IN STD_LOGIC;
    s_axis_tready : OUT STD_LOGIC;
    s_axis_tdata : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    s_axis_tlast : IN STD_LOGIC;
    m_axis_tvalid : OUT STD_LOGIC;
    m_axis_tready : IN STD_LOGIC;
    m_axis_tdata : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    m_axis_tlast : OUT STD_LOGIC;
    axis_prog_full : OUT STD_LOGIC
  );
END COMPONENT;

COMPONENT axi8_fifo_bram
  PORT (
    wr_rst_busy : OUT STD_LOGIC;
    rd_rst_busy : OUT STD_LOGIC;
    m_aclk : IN STD_LOGIC;
    s_aclk : IN STD_LOGIC;
    s_aresetn : IN STD_LOGIC;
    s_axis_tvalid : IN STD_LOGIC;
    s_axis_tready : OUT STD_LOGIC;
    s_axis_tdata : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    s_axis_tlast : IN STD_LOGIC;
    m_axis_tvalid : OUT STD_LOGIC;
    m_axis_tready : IN STD_LOGIC;
    m_axis_tdata : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    m_axis_tlast : OUT STD_LOGIC;
    axis_prog_full : OUT STD_LOGIC
  );
END COMPONENT;

begin
xpm_fifo_gen: if USE_BUILT_IN_FIFO = '0' generate
	axi8_fifo_inst: axi8_fifo_bram
		PORT Map(
			wr_rst_busy 	    => open,
            rd_rst_busy         => open,
            m_aclk              => m_axis_aclk, 
            s_aclk              => s_axis_aclk,
            s_aresetn           => s_axis_aresetn,
            s_axis_tvalid       => s_axis.tvalid,
            s_axis_tready       => s_axis_tready,
            s_axis_tdata        => s_axis.tdata,
            s_axis_tlast        => s_axis.tlast,
            m_axis_tvalid       => m_axis.tvalid,
            m_axis_tready       => m_axis_tready,
            m_axis_tdata        => m_axis.tdata,
            m_axis_tlast        => m_axis.tlast,
            axis_prog_full      => almost_full
        );
--    fifo: xpm_fifo_axis
--        generic map (
--            CLOCKING_MODE => CLOCKING_MODE,
--            FIFO_MEMORY_TYPE => FIFO_MEMORY_TYPE,
--            PACKET_FIFO => PACKET_FIFO,
--            FIFO_DEPTH => DEPTH,
--            TDATA_WIDTH => 8,
--            TID_WIDTH => 1,
--            TDEST_WIDTH => 1,
--            TUSER_WIDTH => 1,
--            ECC_MODE => "no_ecc",
--            RELATED_CLOCKS => RELATED_CLOCKS,
--            USE_ADV_FEATURES => "0008",
--            WR_DATA_COUNT_WIDTH => 1,
--            RD_DATA_COUNT_WIDTH => 1,
--            PROG_FULL_THRESH => DEPTH-2,
--            PROG_EMPTY_THRESH => 5,
--            CDC_SYNC_STAGES => 2
--        )
--        port map (
--            s_aresetn => s_axis_aresetn,
--            m_aclk => m_axis_aclk,
--            s_aclk => s_axis_aclk,
--            s_axis_tvalid => s_axis.tvalid,
--            s_axis_tready => s_axis_tready,
--            s_axis_tdata => s_axis.tdata,
--            s_axis_tstrb => (others => '1'),
--            s_axis_tkeep => (others => '0'),
--            s_axis_tlast => s_axis.tlast,
--            s_axis_tid => (others => '0'),
--            s_axis_tdest => (others => '0'),
--            s_axis_tuser => (others => '0'),
--            m_axis_tvalid => m_axis.tvalid,
--            m_axis_tready => m_axis_tready,
--            m_axis_tdata => m_axis.tdata,
--            m_axis_tstrb => open,
--            m_axis_tkeep => open,
--            m_axis_tlast => m_axis.tlast,
--            m_axis_tid => open,
--            m_axis_tdest => open,
--            m_axis_tuser => open,
--            prog_full_axis => open,
--            wr_data_count_axis => open,
--            almost_full_axis => almost_full,
--            prog_empty_axis => open,
--            rd_data_count_axis => open,
--            almost_empty_axis => open,
--            injectsbiterr_axis => '0',
--            injectdbiterr_axis => '0',
--            sbiterr_axis => open,
--            dbiterr_axis => open
--        );
end generate;
builtin_fifo_gen: if USE_BUILT_IN_FIFO = '1' generate 
    axi8_fifo_inst: axi8_fifo_bif
        PORT Map(
            wr_rst_busy         => open,
            rd_rst_busy         => open,
            m_aclk              => m_axis_aclk, 
            s_aclk              => s_axis_aclk,
            s_aresetn           => s_axis_aresetn,
            s_axis_tvalid       => s_axis.tvalid,
            s_axis_tready       => s_axis_tready,
            s_axis_tdata        => s_axis.tdata,
            s_axis_tlast        => s_axis.tlast,
            m_axis_tvalid       => m_axis.tvalid,
            m_axis_tready       => m_axis_tready,
            m_axis_tdata        => m_axis.tdata,
            m_axis_tlast        => m_axis.tlast,
            axis_prog_full      => almost_full
        );
end generate;
end architecture;
