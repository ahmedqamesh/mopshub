//
// Verilog Module mopshub_lib.canakari_tb
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 12:05:16 01/04/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module canakari_tb ;


// ### Please start your Verilog code here ### 

endmodule
