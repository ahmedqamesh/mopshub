//
// Verilog Module mopshub_reconfig.icap_wrapper
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 10:25:10 05/17/23
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module icap_wrapper ;


// ### Please start your Verilog code here ### 

endmodule
