//
// Verilog Module mopshub_lib.rec_spi_buf_id
//
// Created:
//          by - dcs.dcs (localhost)
//          at - 14:57:24 05/24/22
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module rec_spi_buf_id ;


// ### Please start your Verilog code here ### 

endmodule
