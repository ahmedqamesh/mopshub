//
// Verilog Module mopshub_lib.enc8b10_wrap
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 18:34:27 03/03/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module enc8b10bx ;


// ### Please start your Verilog code here ### 

endmodule
