`resetall
`timescale 1ns/10ps
module can_elink_bridge_SM( 
   // Port Declarations
   input   wire           can_bus_match, 
   input   wire           clk,                 // posedge
   input   wire           end_cnt_dbg, 
   input   wire           end_init,            // Signal from CAN interface block to indicate that initialization process is finished 
   input   wire           end_osc_cnt, 
   input   wire           end_read_can,        // signal from CANopen block to indicate that it has read receive message buffer 
   input   wire           end_read_elink,      // this signal goes high when CANopen block has finshed writing transmit message buffer register 
   input   wire           end_trim_osc, 
   input   wire           end_write_can,       // goes high when can interface block had finished writing canakari transmit registers
   input   wire           end_write_elink,     // Goes high when CANopen block finished reading the received message buffer register 
   input   wire           endwait,             // This signal indicates when message can't be decoded in one of the CANopen objects to go back to known state to receive message
   input   wire           irq_can_rec,         // interrupt signal from canakari to indicate successful read of a new message by one of the 32 buses 
   input   wire           irq_can_tra,         // successful transmission interrupt signal from cankari 
   input   wire           irq_elink_tra,       // interrupt from elink to indicate it has a msg
   input   wire           osc_auto_trim, 
   input   wire    [4:0]  osc_msg_cnt, 
   input   wire           priority_sig, 
   input   wire           reset_irq_rec_done, 
   input   wire           reset_irq_tra_done, 
   input   wire           rst,                 // lowactive
   input   wire           timeoutrst,          // timeout reset in case bridge controller does not respond in a specied amount of time 
   input   wire           timeoutrst_trim,     // timeout reset in case bridge controller does not respond in a specied amount of time 
   output  reg            abort_mes,           // Signals other state machines to come to a known statte 
   output  reg            can_bus_comp, 
   output  reg            can_rec_ack, 
   output  reg            done_trim_osc_all, 
   output  reg            end_can_proc, 
   output  reg            end_trim_bus, 
   output  reg            entimeout,           // enable for timeout reset counter 
   output  reg            entimeout_trim, 
   output  reg            irq_can_ack,         // tto start transmitting CAN message 
   output  reg     [3:0]  mopshub_sm_dbg, 
   output  reg            power_bus_en, 
   output  reg            reset_irq_can,       // reset canakri interrupt 
   output  reg            reset_irq_can_all,   // reset all canakri interrupt 
   output  reg            reset_irq_osc_can, 
   output  reg            reset_irq_rec_can, 
   output  reg            reset_irq_tra_can, 
   output  reg            rst_mops_dbg, 
   output  reg            rst_msg_cnt, 
   output  reg            rst_osc_cnt, 
   output  reg            send_mes_can, 
   output  reg            sign_on_sig,         // Signal to send one time NMT message after bootup
   output  reg            skip_osc_trim, 
   output  reg            start_init,          // to initialize the CAN node (cankari)
   output  reg            start_msg_cnt, 
   output  reg            start_osc_cnt, 
   output  reg            start_read_can,      // to read canakari receive registers
   output  reg            start_read_elink,    // signal to read transmit message buffer register 
   output  reg            start_trim_ack, 
   output  reg            start_trim_osc, 
   output  reg            start_write_can,     // to write transmit registers of canakari 
   output  reg            start_write_elink, 
   output  reg     [5:0]  statedeb
);


// Internal Declarations


// Module Declarations

// State encoding
parameter 
          reset              = 6'd0,
          initialize         = 6'd1,
          waittoact          = 6'd2,
          Abort_current      = 6'd3,
          pass_mes_to_elink  = 6'd4,
          rst_rec_irq_can    = 6'd5,
          write_mes_canakari = 6'd6,
          rst_irq            = 6'd7,
          Wait_tra           = 6'd8,
          read_elink_mes     = 6'd9,
          Wait_for_read      = 6'd10,
          endwaitst          = 6'd11,
          Start              = 6'd12,
          Start_read_new     = 6'd13,
          signon             = 6'd14,
          comp_bus_select    = 6'd15,
          check_rec2         = 6'd16,
          finish_proc        = 6'd17,
          rst_all_irq_can    = 6'd18,
          check_rec1         = 6'd19,
          send_ack           = 6'd20,
          Check_Trim         = 6'd21,
          Wait_for_OSC       = 6'd22,
          s1                 = 6'd23,
          finish_proc1       = 6'd24,
          rst_rec_irq_can1   = 6'd25,
          Rread_Resp         = 6'd26,
          pass_to_elink      = 6'd27,
          Break_Loop         = 6'd28,
          finishtrim         = 6'd29,
          send_ack1          = 6'd30,
          ST_Start_Cnt1      = 6'd31,
          ST_CountRst2       = 6'd32,
          Wait_Resp          = 6'd33,
          rst_irq1           = 6'd34,
          s3                 = 6'd35,
          trim_ack           = 6'd36,
          finish_proc2       = 6'd37,
          RST_MOPS_dbg       = 6'd38,
          s0                 = 6'd39,
          s2                 = 6'd40,
          checkmsg_cnt       = 6'd41,
          Wait_Suc_tra       = 6'd42,
          rst_msg            = 6'd43,
          msg_cnt1           = 6'd44,
          s4                 = 6'd45,
          ST_Skip_Bus        = 6'd46,
          Ack_Receive        = 6'd47;

reg [5:0] current_state, next_state;
// pragma synthesis_off
reg hds_animation_indicator;
// pragma synthesis_on

// Wait State Signals
reg [4:0] csm_timer;
reg [4:0] csm_next_timer;
reg       csm_timeout;
reg       csm_to_Wait_for_read;
reg       csm_to_s0;
reg       csm_to_s4;

//-----------------------------------------------------------------
// Next State Block for machine csm
//-----------------------------------------------------------------
always @(
   can_bus_match, 
   csm_timeout, 
   current_state, 
   end_cnt_dbg, 
   end_init, 
   end_osc_cnt, 
   end_read_can, 
   end_read_elink, 
   end_write_can, 
   end_write_elink, 
   irq_can_rec, 
   irq_can_tra, 
   irq_elink_tra, 
   osc_auto_trim, 
   osc_msg_cnt, 
   priority_sig, 
   reset_irq_rec_done, 
   reset_irq_tra_done, 
   rst
)
begin : next_state_block_proc
   // Default assignments to Wait State entry flags
   csm_to_Wait_for_read = 1'b0;
   csm_to_s0 = 1'b0;
   csm_to_s4 = 1'b0;
   case (current_state) 
      reset: begin
         if (rst == 1) begin
            next_state = Start;
            // pragma synthesis_off
            $hdsNextPath(0,1);
            // pragma synthesis_on
         end
         else begin
            next_state = reset;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      initialize: begin
         if (end_init == 1) begin
            next_state = Wait_for_OSC;
            // pragma synthesis_off
            $hdsNextPath(0,2);
            // pragma synthesis_on
         end
         else begin
            next_state = initialize;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      waittoact: begin
         if (irq_can_rec == 1) begin
            next_state = Wait_for_read;
            csm_to_Wait_for_read = 1'b1;
            // pragma synthesis_off
            $hdsNextPath(0,3);
            // pragma synthesis_on
         end
         else if (irq_elink_tra == 1) begin
            next_state = check_rec1;
            // pragma synthesis_off
            $hdsNextPath(0,4);
            // pragma synthesis_on
         end
         else begin
            next_state = waittoact;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      Abort_current: begin
         next_state = Wait_for_read;
         csm_to_Wait_for_read = 1'b1;
         // pragma synthesis_off
         $hdsNextPath(0,5);
         // pragma synthesis_on
      end
      pass_mes_to_elink: begin
         if (end_write_elink == 1) begin
            next_state = rst_rec_irq_can;
            // pragma synthesis_off
            $hdsNextPath(0,6);
            // pragma synthesis_on
         end
         else begin
            next_state = pass_mes_to_elink;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      rst_rec_irq_can: begin
         if (reset_irq_rec_done ==1) begin
            next_state = finish_proc;
            // pragma synthesis_off
            $hdsNextPath(0,7);
            // pragma synthesis_on
         end
         else begin
            next_state = rst_rec_irq_can;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      write_mes_canakari: begin
         if (end_write_can == 1) begin
            next_state = Wait_tra;
            // pragma synthesis_off
            $hdsNextPath(0,8);
            // pragma synthesis_on
         end
         else begin
            next_state = write_mes_canakari;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      rst_irq: begin
         if (reset_irq_tra_done ==1) begin
            next_state = waittoact;
            // pragma synthesis_off
            $hdsNextPath(0,9);
            // pragma synthesis_on
         end
         else begin
            next_state = rst_irq;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      Wait_tra: begin
         if (irq_can_tra == 1) begin
            next_state = send_ack;
            // pragma synthesis_off
            $hdsNextPath(0,10);
            // pragma synthesis_on
         end
         else begin
            next_state = Wait_tra;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      read_elink_mes: begin
         if (end_read_elink == 1) begin
            next_state = check_rec2;
            // pragma synthesis_off
            $hdsNextPath(0,11);
            // pragma synthesis_on
         end
         else begin
            next_state = read_elink_mes;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      Wait_for_read: begin
         if (csm_timeout) begin
            next_state = Start_read_new;
            // pragma synthesis_off
            $hdsNextPath(0,12);
            // pragma synthesis_on
         end
         else begin
            next_state = Wait_for_read;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      endwaitst: begin
         next_state = rst_all_irq_can;
         // pragma synthesis_off
         $hdsNextPath(0,13);
         // pragma synthesis_on
      end
      Start: begin
         next_state = initialize;
         // pragma synthesis_off
         $hdsNextPath(0,14);
         // pragma synthesis_on
      end
      Start_read_new: begin
         if (end_read_can == 1) begin
            next_state = Ack_Receive;
            // pragma synthesis_off
            $hdsNextPath(0,15);
            // pragma synthesis_on
         end
         else begin
            next_state = Start_read_new;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      signon: begin
         next_state = waittoact;
         // pragma synthesis_off
         $hdsNextPath(0,16);
         // pragma synthesis_on
      end
      comp_bus_select: begin
         if (can_bus_match ==1) begin
            next_state = Wait_for_read;
            csm_to_Wait_for_read = 1'b1;
            // pragma synthesis_off
            $hdsNextPath(0,17);
            // pragma synthesis_on
         end
         else begin
            next_state = read_elink_mes;
            // pragma synthesis_off
            $hdsNextPath(0,18);
            // pragma synthesis_on
         end
      end
      check_rec2: begin
         if (irq_can_rec == 1) begin
            next_state = comp_bus_select;
            // pragma synthesis_off
            $hdsNextPath(0,19);
            // pragma synthesis_on
         end
         else begin
            next_state = write_mes_canakari;
            // pragma synthesis_off
            $hdsNextPath(0,20);
            // pragma synthesis_on
         end
      end
      finish_proc: begin
         next_state = waittoact;
         // pragma synthesis_off
         $hdsNextPath(0,21);
         // pragma synthesis_on
      end
      rst_all_irq_can: begin
         next_state = waittoact;
         // pragma synthesis_off
         $hdsNextPath(0,22);
         // pragma synthesis_on
      end
      check_rec1: begin
         if (priority_sig ==1) begin
            next_state = write_mes_canakari;
            // pragma synthesis_off
            $hdsNextPath(0,23);
            // pragma synthesis_on
         end
         else begin
            next_state = read_elink_mes;
            // pragma synthesis_off
            $hdsNextPath(0,24);
            // pragma synthesis_on
         end
      end
      send_ack: begin
         next_state = rst_irq;
         // pragma synthesis_off
         $hdsNextPath(0,25);
         // pragma synthesis_on
      end
      Check_Trim: begin
         if (osc_auto_trim ==1) begin
            next_state = s3;
            // pragma synthesis_off
            $hdsNextPath(0,26);
            // pragma synthesis_on
         end
         else begin
            next_state = signon;
            // pragma synthesis_off
            $hdsNextPath(0,27);
            // pragma synthesis_on
         end
      end
      Wait_for_OSC: begin
         next_state = Check_Trim;
         // pragma synthesis_off
         $hdsNextPath(0,28);
         // pragma synthesis_on
      end
      s1: begin
         if (end_write_can == 1) begin
            next_state = s2;
            // pragma synthesis_off
            $hdsNextPath(0,29);
            // pragma synthesis_on
         end
         else begin
            next_state = s1;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      finish_proc1: begin
         next_state = finish_proc2;
         // pragma synthesis_off
         $hdsNextPath(0,30);
         // pragma synthesis_on
      end
      rst_rec_irq_can1: begin
         if (reset_irq_rec_done ==1) begin
            next_state = finish_proc1;
            // pragma synthesis_off
            $hdsNextPath(0,31);
            // pragma synthesis_on
         end
         else begin
            next_state = rst_rec_irq_can1;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      Rread_Resp: begin
         if (end_read_can == 1) begin
            next_state = pass_to_elink;
            // pragma synthesis_off
            $hdsNextPath(0,32);
            // pragma synthesis_on
         end
         else begin
            next_state = Rread_Resp;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      pass_to_elink: begin
         if (end_write_elink == 1) begin
            next_state = rst_rec_irq_can1;
            // pragma synthesis_off
            $hdsNextPath(0,33);
            // pragma synthesis_on
         end
         else begin
            next_state = pass_to_elink;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      Break_Loop: begin
         if (end_osc_cnt ==1 |  end_cnt_dbg ==1) begin
            next_state = ST_CountRst2;
            // pragma synthesis_off
            $hdsNextPath(0,34);
            // pragma synthesis_on
         end
         else begin
            next_state = RST_MOPS_dbg;
            // pragma synthesis_off
            $hdsNextPath(0,35);
            // pragma synthesis_on
         end
      end
      finishtrim: begin
         next_state = signon;
         // pragma synthesis_off
         $hdsNextPath(0,36);
         // pragma synthesis_on
      end
      send_ack1: begin
         next_state = rst_irq1;
         // pragma synthesis_off
         $hdsNextPath(0,37);
         // pragma synthesis_on
      end
      ST_Start_Cnt1: begin
         next_state = s3;
         // pragma synthesis_off
         $hdsNextPath(0,38);
         // pragma synthesis_on
      end
      ST_CountRst2: begin
         next_state = s4;
         csm_to_s4 = 1'b1;
         // pragma synthesis_off
         $hdsNextPath(0,39);
         // pragma synthesis_on
      end
      Wait_Resp: begin
         if (irq_can_rec == 1) begin
            next_state = s0;
            csm_to_s0 = 1'b1;
            // pragma synthesis_off
            $hdsNextPath(0,40);
            // pragma synthesis_on
         end
         else begin
            next_state = Wait_Resp;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      rst_irq1: begin
         if (reset_irq_tra_done ==1) begin
            next_state = Wait_Resp;
            // pragma synthesis_off
            $hdsNextPath(0,41);
            // pragma synthesis_on
         end
         else begin
            next_state = rst_irq1;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      s3: begin
         next_state = trim_ack;
         // pragma synthesis_off
         $hdsNextPath(0,42);
         // pragma synthesis_on
      end
      trim_ack: begin
         next_state = s1;
         // pragma synthesis_off
         $hdsNextPath(0,43);
         // pragma synthesis_on
      end
      finish_proc2: begin
         next_state = Break_Loop;
         // pragma synthesis_off
         $hdsNextPath(0,44);
         // pragma synthesis_on
      end
      RST_MOPS_dbg: begin
         next_state = ST_Start_Cnt1;
         // pragma synthesis_off
         $hdsNextPath(0,45);
         // pragma synthesis_on
      end
      s0: begin
         if (csm_timeout) begin
            next_state = Rread_Resp;
            // pragma synthesis_off
            $hdsNextPath(0,46);
            // pragma synthesis_on
         end
         else begin
            next_state = s0;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      s2: begin
         next_state = checkmsg_cnt;
         // pragma synthesis_off
         $hdsNextPath(0,47);
         // pragma synthesis_on
      end
      checkmsg_cnt: begin
         if (osc_msg_cnt ==5'h10) begin
            next_state = rst_msg;
            // pragma synthesis_off
            $hdsNextPath(0,48);
            // pragma synthesis_on
         end
         else begin
            next_state = msg_cnt1;
            // pragma synthesis_off
            $hdsNextPath(0,49);
            // pragma synthesis_on
         end
      end
      Wait_Suc_tra: begin
         if (irq_can_tra ==1) begin
            next_state = send_ack1;
            // pragma synthesis_off
            $hdsNextPath(0,50);
            // pragma synthesis_on
         end
         else begin
            next_state = Wait_Suc_tra;
            // pragma synthesis_off
            $hdsNextPath(0,0);
            // pragma synthesis_on
         end
      end
      rst_msg: begin
         next_state = Wait_Suc_tra;
         // pragma synthesis_off
         $hdsNextPath(0,51);
         // pragma synthesis_on
      end
      msg_cnt1: begin
         next_state = trim_ack;
         // pragma synthesis_off
         $hdsNextPath(0,52);
         // pragma synthesis_on
      end
      s4: begin
         next_state = finishtrim;
         // pragma synthesis_off
         $hdsNextPath(0,53);
         // pragma synthesis_on
      end
      ST_Skip_Bus: begin
         next_state = Break_Loop;
         // pragma synthesis_off
         $hdsNextPath(0,54);
         // pragma synthesis_on
      end
      Ack_Receive: begin
         next_state = pass_mes_to_elink;
         // pragma synthesis_off
         $hdsNextPath(0,55);
         // pragma synthesis_on
      end
      default: begin
         next_state = reset;
         // pragma synthesis_off
         $hdsNextPath(0,0);
         // pragma synthesis_on
      end
   endcase
end // Next State Block

//-----------------------------------------------------------------
// Output Block for machine csm
//-----------------------------------------------------------------
always @(
   current_state
)
begin : output_block_proc
   // Default Assignment
   abort_mes = 0;
   can_bus_comp = 0;
   can_rec_ack = 0;
   done_trim_osc_all = 0;
   end_can_proc = 0;
   end_trim_bus = 0;
   entimeout = 1;
   entimeout_trim = 1;
   irq_can_ack = 0;
   mopshub_sm_dbg = 4'b0;
   power_bus_en = 0;
   reset_irq_can = 0;
   reset_irq_can_all = 0;
   reset_irq_osc_can = 0;
   reset_irq_rec_can = 0;
   reset_irq_tra_can = 0;
   rst_mops_dbg = 0;
   rst_msg_cnt = 0;
   rst_osc_cnt = 0;
   send_mes_can = 0;
   sign_on_sig = 0;
   skip_osc_trim = 0;
   start_init = 0;
   start_msg_cnt = 0;
   start_osc_cnt = 0;
   start_read_can = 0;
   start_read_elink = 0;
   start_trim_ack = 0;
   start_trim_osc = 0;
   start_write_can = 0;
   start_write_elink = 0;

   // Combined Actions
   case (current_state) 
      reset: begin
         abort_mes = 1 ;
         reset_irq_can = 0 ;
         reset_irq_can_all = 0 ;
         send_mes_can = 0 ;  
         start_read_can = 0 ;
         start_read_elink = 0 ;
         start_write_can = 0 ;
         start_write_elink = 0 ;
         start_init = 0 ;
         sign_on_sig = 0;
         entimeout = 0 ;
         entimeout_trim = 0;
         skip_osc_trim = 0;
         can_rec_ack =0;
      end
      initialize: begin
         start_init = 1 ;
         entimeout = 0 ;
         entimeout_trim =0;
      end
      waittoact: begin
         entimeout = 0 ;
         entimeout_trim = 0;
         mopshub_sm_dbg =4'b001;
      end
      Abort_current: begin
         abort_mes = 1 ;
      end
      pass_mes_to_elink: begin
         start_write_elink = 1;
         mopshub_sm_dbg =4'b011;
      end
      rst_rec_irq_can: begin
         reset_irq_can = 1 ;
         reset_irq_rec_can = 1 ;
         mopshub_sm_dbg =4'b100;
      end
      write_mes_canakari: begin
         start_write_can = 1 ;
         mopshub_sm_dbg =4'b111;
      end
      rst_irq: begin
         reset_irq_can = 1 ;
         reset_irq_tra_can = 1 ;
         mopshub_sm_dbg =4'b1010;
      end
      Wait_tra: begin
         send_mes_can =1;
         mopshub_sm_dbg =4'b1000;
      end
      read_elink_mes: begin
         start_read_elink = 1 ;
      end
      Start_read_new: begin
         start_read_can = 1 ;
         mopshub_sm_dbg =4'b010;
      end
      signon: begin
         sign_on_sig = 1 ;
      end
      comp_bus_select: begin
         can_bus_comp =1;
      end
      finish_proc: begin
         end_can_proc = 1;
         mopshub_sm_dbg =4'b101;
      end
      rst_all_irq_can: begin
         reset_irq_can_all = 1 ;
      end
      check_rec1: begin
         mopshub_sm_dbg =4'b110;
      end
      send_ack: begin
         irq_can_ack = 1 ;
         mopshub_sm_dbg =4'b1001;
      end
      s1: begin
         start_trim_osc =1;
      end
      finish_proc1: begin
         end_can_proc = 1;
      end
      rst_rec_irq_can1: begin
         reset_irq_can = 1 ;
         reset_irq_rec_can = 1 ;
      end
      Rread_Resp: begin
         start_read_can = 1 ;
      end
      pass_to_elink: begin
         start_write_elink = 1;
      end
      finishtrim: begin
         done_trim_osc_all =1;
      end
      send_ack1: begin
         irq_can_ack = 1 ;
      end
      ST_Start_Cnt1: begin
         start_osc_cnt =1;
      end
      ST_CountRst2: begin
         rst_osc_cnt =1;
      end
      Wait_Resp: begin
         entimeout =0;
      end
      rst_irq1: begin
         reset_irq_can = 1 ;
         reset_irq_osc_can = 1 ;
      end
      s3: begin
         power_bus_en =1;
      end
      trim_ack: begin
         start_trim_ack =1;
      end
      finish_proc2: begin
         end_trim_bus =1;
      end
      RST_MOPS_dbg: begin
         rst_mops_dbg =1;
      end
      s2: begin
         send_mes_can =1;
      end
      Wait_Suc_tra: begin
         entimeout =0;
      end
      rst_msg: begin
         rst_msg_cnt  = 1;
      end
      msg_cnt1: begin
         start_msg_cnt  = 1;
      end
      ST_Skip_Bus: begin
         entimeout_trim =0;
         skip_osc_trim = 1;
      end
      Ack_Receive: begin
         can_rec_ack = 1;
      end
   endcase
end // Output Block

//-----------------------------------------------------------------
// Clocked Block for machine csm
//-----------------------------------------------------------------
always @(
   posedge clk, 
   negedge rst
) 
begin : clocked_block_proc
   if (!rst) begin
      current_state <= reset;
      csm_timer <= 5'd0;
   end
   else 
   begin
      if (endwait) begin
         current_state <= reset;
         csm_timer <= 5'd0;
      end
      else if (timeoutrst) begin
         current_state <= endwaitst;
         csm_timer <= 5'd0;
      end
      else if (timeoutrst_trim) begin
         current_state <= ST_Skip_Bus;
         csm_timer <= 5'd0;
      end
      else 
      begin
         current_state <= next_state;
         csm_timer <= csm_next_timer;
         // pragma synthesis_off
         $hdsClock(0);
         // pragma synthesis_on
      end
   end
end // Clocked Block

//-----------------------------------------------------------------
// Wait state logic for machine csm
//-----------------------------------------------------------------
always @(
   csm_timer,
   csm_to_Wait_for_read,
   csm_to_s0,
   csm_to_s4
)
begin : csm_wait_block_proc
   csm_timeout = (csm_timer == 5'd0);
   if (csm_to_Wait_for_read == 1'b1) begin
      csm_next_timer = 5'd19;  //no cycles(20)-1=19
   end
   else if (csm_to_s0 == 1'b1) begin
      csm_next_timer = 5'd19;  //no cycles(20)-1=19
   end
   else if (csm_to_s4 == 1'b1) begin
      csm_next_timer = 5'd19;  //no cycles(20)-1=19
   end
   else begin
      csm_next_timer = (csm_timeout)? 5'd0: (csm_timer - 5'd1);
   end
end // Wait State Block
// State-As-Output assignment
always @(current_state)
statedeb = current_state;

endmodule // can_elink_bridge_SM
