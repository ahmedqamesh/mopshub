`resetall
`timescale 1ns/10ps
module tb_mopshub_top();
  wire              clk ;//= 1'b0;
  wire             clk_40;
  wire             clk_80;
  reg             rst   = 1'b1;
  wire            rst_mops_dbg;
  reg             sel_bus = 1'b0;
  reg     [4:0]   can_tra_select_dbg =5'd1;
  wire            sign_on_sig;
  reg             start_data_gen= 1'b0;
  wire            start_init;
  wire            end_init;
  string          info_debug_sig;     
  //tbSM signals  
  wire    [75:0]  bus_dec_data;
  wire    [7:0]   bus_id;
  int             adc_ch;
  
  //Automated trimming signals
  reg             osc_auto_trim =1'b0; ////Active high. Enable /disable automated trimming. If disabled then take care of ftrim_pads_reg
  wire            trim_sig_start;
  wire            trim_sig_end;
  wire            trim_sig_done;
  
  reg             osc_auto_trim_mopshub =1'b0;
  wire            ready_osc;
  wire            start_trim_osc;
  wire            end_trim_bus;
  wire            done_trim_osc;
  
  wire            power_bus_en;
  wire    [4:0]   power_bus_cnt;
  
  wire            sign_in_start;
  wire            sign_in_end;
  reg             test_rx = 1'b0;
  wire            test_rx_start;
  wire            test_rx_end;
  
  reg             test_tx = 1'b0;
  wire            test_tx_start;
  wire            test_tx_end;
  
  // MOPSHUB signals
  wire    [75:0]  data_rec_uplink;
  wire    [75:0]  data_tra_emulator_out;
  wire    [4:0]   can_rec_select;
  wire    [75:0]  data_tra_downlink;
  wire    [4:0]  can_tra_select;
  wire    [75:0] data_rec_emulator_in;
  wire            irq_elink_tra;
  wire            irq_elink_rec;
  
  // Generator signals 
  wire            rx0;
  wire            rx1;
  wire            rx2;
  wire            rx3;
  wire            rx4;
  wire            rx5;
  wire            rx6;
  wire            rx7;
  
  wire            tx0;
  wire            tx1;
  wire            tx2;
  wire            tx3;
  wire            tx4;
  wire            tx5;
  wire            tx6;
  wire            tx7;
  //wire [1:0] tx_mopshub_2bit; 
  wire       tx_mopshub_1bit; 
  //wire [1:0] rx_mopshub_2bit; 
  wire       rx_mopshub_1bit;
  
  //Internal assignments  
  assign can_tra_select   = mopshub0.can_tra_select;
  assign can_rec_select   = mopshub0.can_rec_select;
  assign data_rec_uplink  = mopshub0.data_rec_uplink;
  assign data_tra_downlink  = mopshub0.data_tra_downlink;
  assign done_trim_osc    = mopshub0.done_trim_osc;
  assign start_init       = mopshub0.start_init;
  assign end_init         = mopshub0.end_init;
  assign rst_mops_dbg     = mopshub0.rst_mops_dbg;
  assign sign_on_sig      = mopshub0.sign_on_sig;
  assign end_trim_bus     = mopshub0.end_trim_bus;
  assign start_trim_osc   = mopshub0.start_trim_ack;
  assign power_bus_en     = mopshub0.power_bus_en;
  assign power_bus_cnt    = mopshub0.power_bus_cnt;  
  assign irq_elink_tra    = mopshub0.irq_elink_tra;
  assign irq_elink_rec    = mopshub0.irq_elink_rec;
  assign data_tra_emulator_out  = data_generator0.data_tra_76bit_reg;
  assign data_rec_emulator_in   = data_generator0.data_rec_76bit_reg;
  assign ready_osc              = data_generator0.ready_osc;
  
  
  mopshub_top#(
  .n_buses (5'b111),
  .seialize_data_stream(1),
  .generate_mopshub(1'b1))mopshub0(
  .clk(clk_40),
  .clk_80(clk_80),
  .reset(!rst),  
  .osc_auto_trim_mopshub(osc_auto_trim_mopshub),                     
  .end_cnt_dbg(1'b0),      
  //.tx_elink2bit(tx_mopshub_2bit),
  .tx_elink1bit(tx_mopshub_1bit),
  .rx_elink1bit(rx_mopshub_1bit),
  // .rx_elink2bit(rx_mopshub_2bit),        
  .rx0(rx0),        
  .rx1(rx1),        
  .rx2(rx2),        
  .rx3(rx3),        
  .rx4(rx4),        
  .rx5(rx5),        
  .rx6(rx6),        
  .rx7(rx7),
  .tx0(tx0),              
  .tx1(tx1),
  .tx2(tx2),
  .tx3(tx3),
  .tx4(tx4),
  .tx5(tx5),
  .tx6(tx6),
  .tx7(tx7));
  
  data_generator#(
  .n_buses (5'b111),
  .seialize_data_stream(1),
  .generate_mopshub(1'b1))data_generator0(
  .clk(clk_40),
  .clk_80(clk_80),
  .rst(rst),
  .ext_rst_mops(rst_mops_dbg),
  .ext_trim_mops(osc_auto_trim_mopshub),
  .loop_en(1'b0),
  //Start SM
  .start_data_gen(start_data_gen),
  //OScillation Triming Signals
  .osc_auto_trim(osc_auto_trim),
  .trim_sig_start(trim_sig_start),
  .trim_sig_end (trim_sig_end),
  .trim_sig_done(trim_sig_done),
  .sign_in_start(sign_in_start), 
  .sign_in_end(sign_in_end),
  //Read ADC channels from MOPS and send it to MOPSHUB rx
  .test_rx(test_rx),
  .test_tx(test_tx),
  .test_tx_end(test_tx_end),
  .test_rx_start(test_rx_start),
  .test_rx_end(test_rx_end),
  .test_tx_start(test_tx_start),
  .respmsg(respmsg),
  .reqmsg(reqmsg),
  .adc_ch(adc_ch),  
  // Acknowledgement bit from the MOPSHUB
  //Decoder Signals [Listen always to the bus ]
  .bus_dec_data(bus_dec_data),
  .power_bus_cnt(power_bus_cnt),
  //read data from Elink and send it to the bus
  .sel_bus(sel_bus),
  .bus_cnt(can_tra_select_dbg),// test Bus 0
  .test_mopshub_core(1'b0),
  .osc_auto_trim_mopshub(osc_auto_trim_mopshub),
  .can_rec_select(can_rec_select),
  .bus_id(bus_id),
  .buffer_en(),
  .test_elink_data_done(),
  .start_write_emulator(),
  .start_read_elink(),
  .end_read_elink(),
  //print activity
  .start_init(start_init),   
  .end_init(end_init),
  .can_tra_select(can_tra_select),
  .data_rec_uplink(data_rec_uplink), 
  .data_tra_downlink(data_tra_downlink), 
  .end_trim_bus(end_trim_bus),
  .start_trim_osc(start_trim_osc),
  //Elin.kSignals
  .tx_elink1bit(rx_mopshub_1bit),
  // .tx_elink2bit(rx_mopshub_2bit),
  .rx_elink1bit(tx_mopshub_1bit),
  // .rx_elink2bit(tx_mopshub_2bit),
  //RX-TX signals
  .rx0(rx0),        
  .rx1(rx1),        
  .rx2(rx2),        
  .rx3(rx3),        
  .rx4(rx4),        
  .rx5(rx5),        
  .rx6(rx6),        
  .rx7(rx7),
  .tx0(tx0),              
  .tx1(tx1),
  .tx2(tx2),
  .tx3(tx3),
  .tx4(tx4),
  .tx5(tx5),
  .tx6(tx6),
  .tx7(tx7));
  
  
  //Clock Generators and Dividers
  clock_generator #(
  .freq(40))
  clock_generator0( 
  .clk  (clk), 
  .enable (1'b1)
  ); 
  
  clock_divider #(28'd4)
  clock_divider4( 
  .clock_in  (clk), 
  .clock_out (clk_40)
  ); 
  
  
  clock_divider #(28'd2)
  clock_divider2( 
  .clock_in  (clk), 
  .clock_out (clk_80)
  ); 
  /////******* Reset Generator task--low active ****/////
  initial 
  begin
    rst = 1'b0;
    #10
    rst = 1'b1;
  end
  always@(posedge sign_on_sig)
  begin
    #1500
    start_data_gen = 1'b1;
    #100
    start_data_gen = 1'b0;
  end  
  /////*******Start Full SM for Data Generation ****/////
  always@(posedge clk_40)
  begin  
    if(trim_sig_done ==1 ||done_trim_osc ==1)
    begin
      osc_auto_trim =1'b0;
      osc_auto_trim_mopshub = 1'b0;
    end
    if(sign_on_sig ==1)//start Rx test
    begin
      start_data_gen =1'b0;
      test_tx =1'b1;
    end
    if(test_rx_end ==1)//Done Rx test
    begin
      test_rx =1'b0;
      test_tx =1'b1; 
    end
    if (test_tx_end ==1)//Done Tx test
    test_tx =1'b0;
  end
  
  /////******* prints bus activity ******///
  always@(posedge clk_40)
  if (!rst)
  begin
    info_debug_sig = "<:RESET>";
  end
  else 
  begin
    if(start_init)
    begin 
      info_debug_sig = "<:initialization:>";
    end     
    /////*********************************Oscillator Trimming*********************************///// 
    if(start_trim_osc)
    begin 
      info_debug_sig = {"<:Oscillator Trimming [BUS ID ",$sformatf("%h",power_bus_cnt)," ]:>"};
    end
    if(trim_sig_start)
    begin 
      info_debug_sig = {"<:Oscillator Trimming [BUS ID ",$sformatf("%h",bus_id)," ]:>"};
    end       
    /////*********************************  RX Test    *********************************///// 
    if(test_rx_start)
    begin 
      info_debug_sig = $sformatf("<:RX signals   [BUS ID %d ]  :>",bus_id);
    end 
    /////*********************************  TX Test    *********************************/////     
    if (test_tx_start)
    begin 
      info_debug_sig = $sformatf("<:TX signals  [BUS ID %d ]  :>",bus_id);
    end     
    if(test_tx_end || test_rx_end ||end_init||(end_trim_bus||trim_sig_end))
    begin 
      info_debug_sig = {""};
    end    
  end
endmodule 
