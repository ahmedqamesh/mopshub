//
// Verilog Module mopshub_lib.testbench_tester
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 13:24:46 01/07/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module testbench_tester ;


// ### Please start your Verilog code here ### 

endmodule
