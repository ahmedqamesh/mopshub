//
// Verilog Module mopshub_lib.buffer_tra_spi_data
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 12:04:40 01/27/22
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module buffer_tra_spi_data( 
   // Port Declarations
   input   wire            clk, 
   input   wire    [31:0]  data_tra_in,   // input data from the SCB or Object Dictionary side
   input   wire            buffer_en,     // enable signal
   input   wire            rst, 
   output  wire    [7:0]   spi_id,
   output  wire    [7:0]   spi_reg,
   output  wire    [7:0]   spi_select,
   output  wire    [7:0]   data_tra_out   // Output data to be written on the CAN bus
);

// Internal Declarations
reg [7:0] data_tra_reg   = 8'd0 ;
reg [7:0] spi_id_reg     = 8'd0;
reg [7:0] spi_reg_reg    = 8'd0;
reg [7:0] spi_select_reg = 8'd0;


always@(posedge clk)
begin 
 if(!rst) spi_id_reg <= 8'd0;
 else
  if(buffer_en) spi_id_reg <= data_tra_in[31:24];
  else  spi_id_reg <= spi_id_reg;
end 

always@(posedge clk)
begin 
 if(!rst) spi_select_reg <= 8'd0;
 else
  if(buffer_en) spi_select_reg <= data_tra_in[23:16];
  else  spi_select_reg <= spi_select_reg;
end 

always@(posedge clk)
begin 
 if(!rst) spi_reg_reg <= 8'd0;
 else
  if(buffer_en) spi_reg_reg <= data_tra_in[15:8] ;
  else  spi_reg_reg <= spi_reg_reg;
end 



always@(posedge clk)
begin 
 if(!rst) data_tra_reg <= 8'd0;
 else
  if(buffer_en) data_tra_reg <= data_tra_in[7:0];
  else  data_tra_reg <= data_tra_reg;
end 

assign data_tra_out = data_tra_reg;
assign spi_id = spi_id_reg;
assign spi_reg = spi_reg_reg;
assign spi_select = spi_select_reg;
endmodule
