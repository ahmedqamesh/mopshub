//
// Verilog Module mopshub_lib.canakari_bus_debugger
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 17:23:21 07/21/21
//
// using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
//

`resetall
`timescale 1ns/10ps
module canakari_bus_debugger ;


// ### Please start your Verilog code here ### 

endmodule
