//
// Verilog Module mopshub_lib.elinkRXfifo_wrap
//
// Created:
//          by - dcs.dcs (chipdev2.physik.uni-wuppertal.de)
//          at - 19:45:10 04/02/21
//
// using Mentor Graphics HDL Designer(TM) 2018.1 (Build 12)
//

`resetall
`timescale 1ns/10ps
module elinkRXfifo_wrap(
       // -----------------------------
       // ------ General Interface ---- 
        input   wire           bitClk, 
        input   wire           rst, 
        input   wire           inhibit, 
        input   wire           flush_fifo, 
       // -----------------------------
       // ---- EPROC_IN2 Interface ----
        input   wire    [9:0]  din, 
        input   wire           din_rdy, 
        input   wire           swap_inputbits,
       // ----------------------------
       // --- User Logic Interface ---
        input   wire           rd_clk_elink, 
        input   wire           rd_en_elink, 
        output  wire           empty_elink, 
        output  wire           full_elink, 
        output   wire    [9:0]  dout_elink 
);
// ### Please start your Verilog code here ### 

endmodule
